
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"04",x"07",x"03"),
     1 => (x"74",x"20",x"00",x"00"),
     2 => (x"78",x"7c",x"54",x"54"),
     3 => (x"7f",x"7f",x"00",x"00"),
     4 => (x"38",x"7c",x"44",x"44"),
     5 => (x"7c",x"38",x"00",x"00"),
     6 => (x"00",x"44",x"44",x"44"),
     7 => (x"7c",x"38",x"00",x"00"),
     8 => (x"7f",x"7f",x"44",x"44"),
     9 => (x"7c",x"38",x"00",x"00"),
    10 => (x"18",x"5c",x"54",x"54"),
    11 => (x"7e",x"04",x"00",x"00"),
    12 => (x"00",x"05",x"05",x"7f"),
    13 => (x"bc",x"18",x"00",x"00"),
    14 => (x"7c",x"fc",x"a4",x"a4"),
    15 => (x"7f",x"7f",x"00",x"00"),
    16 => (x"78",x"7c",x"04",x"04"),
    17 => (x"00",x"00",x"00",x"00"),
    18 => (x"00",x"40",x"7d",x"3d"),
    19 => (x"80",x"80",x"00",x"00"),
    20 => (x"00",x"7d",x"fd",x"80"),
    21 => (x"7f",x"7f",x"00",x"00"),
    22 => (x"44",x"6c",x"38",x"10"),
    23 => (x"00",x"00",x"00",x"00"),
    24 => (x"00",x"40",x"7f",x"3f"),
    25 => (x"0c",x"7c",x"7c",x"00"),
    26 => (x"78",x"7c",x"0c",x"18"),
    27 => (x"7c",x"7c",x"00",x"00"),
    28 => (x"78",x"7c",x"04",x"04"),
    29 => (x"7c",x"38",x"00",x"00"),
    30 => (x"38",x"7c",x"44",x"44"),
    31 => (x"fc",x"fc",x"00",x"00"),
    32 => (x"18",x"3c",x"24",x"24"),
    33 => (x"3c",x"18",x"00",x"00"),
    34 => (x"fc",x"fc",x"24",x"24"),
    35 => (x"7c",x"7c",x"00",x"00"),
    36 => (x"08",x"0c",x"04",x"04"),
    37 => (x"5c",x"48",x"00",x"00"),
    38 => (x"20",x"74",x"54",x"54"),
    39 => (x"3f",x"04",x"00",x"00"),
    40 => (x"00",x"44",x"44",x"7f"),
    41 => (x"7c",x"3c",x"00",x"00"),
    42 => (x"7c",x"7c",x"40",x"40"),
    43 => (x"3c",x"1c",x"00",x"00"),
    44 => (x"1c",x"3c",x"60",x"60"),
    45 => (x"60",x"7c",x"3c",x"00"),
    46 => (x"3c",x"7c",x"60",x"30"),
    47 => (x"38",x"6c",x"44",x"00"),
    48 => (x"44",x"6c",x"38",x"10"),
    49 => (x"bc",x"1c",x"00",x"00"),
    50 => (x"1c",x"3c",x"60",x"e0"),
    51 => (x"64",x"44",x"00",x"00"),
    52 => (x"44",x"4c",x"5c",x"74"),
    53 => (x"08",x"08",x"00",x"00"),
    54 => (x"41",x"41",x"77",x"3e"),
    55 => (x"00",x"00",x"00",x"00"),
    56 => (x"00",x"00",x"7f",x"7f"),
    57 => (x"41",x"41",x"00",x"00"),
    58 => (x"08",x"08",x"3e",x"77"),
    59 => (x"01",x"01",x"02",x"00"),
    60 => (x"01",x"02",x"02",x"03"),
    61 => (x"7f",x"7f",x"7f",x"00"),
    62 => (x"7f",x"7f",x"7f",x"7f"),
    63 => (x"1c",x"08",x"08",x"00"),
    64 => (x"7f",x"3e",x"3e",x"1c"),
    65 => (x"3e",x"7f",x"7f",x"7f"),
    66 => (x"08",x"1c",x"1c",x"3e"),
    67 => (x"18",x"10",x"00",x"08"),
    68 => (x"10",x"18",x"7c",x"7c"),
    69 => (x"30",x"10",x"00",x"00"),
    70 => (x"10",x"30",x"7c",x"7c"),
    71 => (x"60",x"30",x"10",x"00"),
    72 => (x"06",x"1e",x"78",x"60"),
    73 => (x"3c",x"66",x"42",x"00"),
    74 => (x"42",x"66",x"3c",x"18"),
    75 => (x"6a",x"38",x"78",x"00"),
    76 => (x"38",x"6c",x"c6",x"c2"),
    77 => (x"00",x"00",x"60",x"00"),
    78 => (x"60",x"00",x"00",x"60"),
    79 => (x"5b",x"5e",x"0e",x"00"),
    80 => (x"1e",x"0e",x"5d",x"5c"),
    81 => (x"ee",x"c2",x"4c",x"71"),
    82 => (x"c0",x"4d",x"bf",x"d5"),
    83 => (x"74",x"1e",x"c0",x"4b"),
    84 => (x"87",x"c7",x"02",x"ab"),
    85 => (x"c0",x"48",x"a6",x"c4"),
    86 => (x"c4",x"87",x"c5",x"78"),
    87 => (x"78",x"c1",x"48",x"a6"),
    88 => (x"73",x"1e",x"66",x"c4"),
    89 => (x"87",x"df",x"ee",x"49"),
    90 => (x"e0",x"c0",x"86",x"c8"),
    91 => (x"87",x"ef",x"ef",x"49"),
    92 => (x"6a",x"4a",x"a5",x"c4"),
    93 => (x"87",x"f0",x"f0",x"49"),
    94 => (x"cb",x"87",x"c6",x"f1"),
    95 => (x"c8",x"83",x"c1",x"85"),
    96 => (x"ff",x"04",x"ab",x"b7"),
    97 => (x"26",x"26",x"87",x"c7"),
    98 => (x"26",x"4c",x"26",x"4d"),
    99 => (x"1e",x"4f",x"26",x"4b"),
   100 => (x"ee",x"c2",x"4a",x"71"),
   101 => (x"ee",x"c2",x"5a",x"d9"),
   102 => (x"78",x"c7",x"48",x"d9"),
   103 => (x"87",x"dd",x"fe",x"49"),
   104 => (x"73",x"1e",x"4f",x"26"),
   105 => (x"c0",x"4a",x"71",x"1e"),
   106 => (x"d3",x"03",x"aa",x"b7"),
   107 => (x"e0",x"d4",x"c2",x"87"),
   108 => (x"87",x"c4",x"05",x"bf"),
   109 => (x"87",x"c2",x"4b",x"c1"),
   110 => (x"d4",x"c2",x"4b",x"c0"),
   111 => (x"87",x"c4",x"5b",x"e4"),
   112 => (x"5a",x"e4",x"d4",x"c2"),
   113 => (x"bf",x"e0",x"d4",x"c2"),
   114 => (x"c1",x"9a",x"c1",x"4a"),
   115 => (x"ec",x"49",x"a2",x"c0"),
   116 => (x"48",x"fc",x"87",x"e8"),
   117 => (x"bf",x"e0",x"d4",x"c2"),
   118 => (x"87",x"ef",x"fe",x"78"),
   119 => (x"c4",x"4a",x"71",x"1e"),
   120 => (x"49",x"72",x"1e",x"66"),
   121 => (x"26",x"87",x"ee",x"ea"),
   122 => (x"71",x"1e",x"4f",x"26"),
   123 => (x"48",x"d4",x"ff",x"4a"),
   124 => (x"ff",x"78",x"ff",x"c3"),
   125 => (x"e1",x"c0",x"48",x"d0"),
   126 => (x"48",x"d4",x"ff",x"78"),
   127 => (x"49",x"72",x"78",x"c1"),
   128 => (x"78",x"71",x"31",x"c4"),
   129 => (x"c0",x"48",x"d0",x"ff"),
   130 => (x"4f",x"26",x"78",x"e0"),
   131 => (x"e0",x"d4",x"c2",x"1e"),
   132 => (x"d1",x"e6",x"49",x"bf"),
   133 => (x"cd",x"ee",x"c2",x"87"),
   134 => (x"78",x"bf",x"e8",x"48"),
   135 => (x"48",x"c9",x"ee",x"c2"),
   136 => (x"c2",x"78",x"bf",x"ec"),
   137 => (x"4a",x"bf",x"cd",x"ee"),
   138 => (x"99",x"ff",x"c3",x"49"),
   139 => (x"72",x"2a",x"b7",x"c8"),
   140 => (x"c2",x"b0",x"71",x"48"),
   141 => (x"26",x"58",x"d5",x"ee"),
   142 => (x"5b",x"5e",x"0e",x"4f"),
   143 => (x"71",x"0e",x"5d",x"5c"),
   144 => (x"87",x"c8",x"ff",x"4b"),
   145 => (x"48",x"c8",x"ee",x"c2"),
   146 => (x"49",x"73",x"50",x"c0"),
   147 => (x"70",x"87",x"f7",x"e5"),
   148 => (x"9c",x"c2",x"4c",x"49"),
   149 => (x"cb",x"49",x"ee",x"cb"),
   150 => (x"49",x"70",x"87",x"ce"),
   151 => (x"c8",x"ee",x"c2",x"4d"),
   152 => (x"c1",x"05",x"bf",x"97"),
   153 => (x"66",x"d0",x"87",x"e2"),
   154 => (x"d1",x"ee",x"c2",x"49"),
   155 => (x"d6",x"05",x"99",x"bf"),
   156 => (x"49",x"66",x"d4",x"87"),
   157 => (x"bf",x"c9",x"ee",x"c2"),
   158 => (x"87",x"cb",x"05",x"99"),
   159 => (x"c5",x"e5",x"49",x"73"),
   160 => (x"02",x"98",x"70",x"87"),
   161 => (x"c1",x"87",x"c1",x"c1"),
   162 => (x"87",x"c0",x"fe",x"4c"),
   163 => (x"e3",x"ca",x"49",x"75"),
   164 => (x"02",x"98",x"70",x"87"),
   165 => (x"ee",x"c2",x"87",x"c6"),
   166 => (x"50",x"c1",x"48",x"c8"),
   167 => (x"97",x"c8",x"ee",x"c2"),
   168 => (x"e3",x"c0",x"05",x"bf"),
   169 => (x"d1",x"ee",x"c2",x"87"),
   170 => (x"66",x"d0",x"49",x"bf"),
   171 => (x"d6",x"ff",x"05",x"99"),
   172 => (x"c9",x"ee",x"c2",x"87"),
   173 => (x"66",x"d4",x"49",x"bf"),
   174 => (x"ca",x"ff",x"05",x"99"),
   175 => (x"e4",x"49",x"73",x"87"),
   176 => (x"98",x"70",x"87",x"c4"),
   177 => (x"87",x"ff",x"fe",x"05"),
   178 => (x"fa",x"fa",x"48",x"74"),
   179 => (x"5b",x"5e",x"0e",x"87"),
   180 => (x"f8",x"0e",x"5d",x"5c"),
   181 => (x"4c",x"4d",x"c0",x"86"),
   182 => (x"c4",x"7e",x"bf",x"ec"),
   183 => (x"ee",x"c2",x"48",x"a6"),
   184 => (x"c1",x"78",x"bf",x"d5"),
   185 => (x"c7",x"1e",x"c0",x"1e"),
   186 => (x"87",x"cd",x"fd",x"49"),
   187 => (x"98",x"70",x"86",x"c8"),
   188 => (x"ff",x"87",x"cd",x"02"),
   189 => (x"87",x"ea",x"fa",x"49"),
   190 => (x"e3",x"49",x"da",x"c1"),
   191 => (x"4d",x"c1",x"87",x"c8"),
   192 => (x"97",x"c8",x"ee",x"c2"),
   193 => (x"87",x"cf",x"02",x"bf"),
   194 => (x"bf",x"d8",x"d4",x"c2"),
   195 => (x"c2",x"b9",x"c1",x"49"),
   196 => (x"71",x"59",x"dc",x"d4"),
   197 => (x"c2",x"87",x"d3",x"fb"),
   198 => (x"4b",x"bf",x"cd",x"ee"),
   199 => (x"bf",x"e0",x"d4",x"c2"),
   200 => (x"87",x"e9",x"c0",x"05"),
   201 => (x"e2",x"49",x"fd",x"c3"),
   202 => (x"fa",x"c3",x"87",x"dc"),
   203 => (x"87",x"d6",x"e2",x"49"),
   204 => (x"ff",x"c3",x"49",x"73"),
   205 => (x"c0",x"1e",x"71",x"99"),
   206 => (x"87",x"e0",x"fa",x"49"),
   207 => (x"b7",x"c8",x"49",x"73"),
   208 => (x"c1",x"1e",x"71",x"29"),
   209 => (x"87",x"d4",x"fa",x"49"),
   210 => (x"f5",x"c5",x"86",x"c8"),
   211 => (x"d1",x"ee",x"c2",x"87"),
   212 => (x"02",x"9b",x"4b",x"bf"),
   213 => (x"d4",x"c2",x"87",x"dd"),
   214 => (x"c7",x"49",x"bf",x"dc"),
   215 => (x"98",x"70",x"87",x"d6"),
   216 => (x"c0",x"87",x"c4",x"05"),
   217 => (x"c2",x"87",x"d2",x"4b"),
   218 => (x"fb",x"c6",x"49",x"e0"),
   219 => (x"e0",x"d4",x"c2",x"87"),
   220 => (x"c2",x"87",x"c6",x"58"),
   221 => (x"c0",x"48",x"dc",x"d4"),
   222 => (x"c2",x"49",x"73",x"78"),
   223 => (x"87",x"cd",x"05",x"99"),
   224 => (x"e1",x"49",x"eb",x"c3"),
   225 => (x"49",x"70",x"87",x"c0"),
   226 => (x"c2",x"02",x"99",x"c2"),
   227 => (x"73",x"4c",x"fb",x"87"),
   228 => (x"05",x"99",x"c1",x"49"),
   229 => (x"f4",x"c3",x"87",x"cd"),
   230 => (x"87",x"ea",x"e0",x"49"),
   231 => (x"99",x"c2",x"49",x"70"),
   232 => (x"fa",x"87",x"c2",x"02"),
   233 => (x"c8",x"49",x"73",x"4c"),
   234 => (x"87",x"cd",x"05",x"99"),
   235 => (x"e0",x"49",x"f5",x"c3"),
   236 => (x"49",x"70",x"87",x"d4"),
   237 => (x"d5",x"02",x"99",x"c2"),
   238 => (x"d9",x"ee",x"c2",x"87"),
   239 => (x"87",x"ca",x"02",x"bf"),
   240 => (x"c2",x"88",x"c1",x"48"),
   241 => (x"c0",x"58",x"dd",x"ee"),
   242 => (x"4c",x"ff",x"87",x"c2"),
   243 => (x"49",x"73",x"4d",x"c1"),
   244 => (x"ce",x"05",x"99",x"c4"),
   245 => (x"49",x"f2",x"c3",x"87"),
   246 => (x"87",x"ea",x"df",x"ff"),
   247 => (x"99",x"c2",x"49",x"70"),
   248 => (x"c2",x"87",x"dc",x"02"),
   249 => (x"7e",x"bf",x"d9",x"ee"),
   250 => (x"a8",x"b7",x"c7",x"48"),
   251 => (x"87",x"cb",x"c0",x"03"),
   252 => (x"80",x"c1",x"48",x"6e"),
   253 => (x"58",x"dd",x"ee",x"c2"),
   254 => (x"fe",x"87",x"c2",x"c0"),
   255 => (x"c3",x"4d",x"c1",x"4c"),
   256 => (x"df",x"ff",x"49",x"fd"),
   257 => (x"49",x"70",x"87",x"c0"),
   258 => (x"d5",x"02",x"99",x"c2"),
   259 => (x"d9",x"ee",x"c2",x"87"),
   260 => (x"c9",x"c0",x"02",x"bf"),
   261 => (x"d9",x"ee",x"c2",x"87"),
   262 => (x"c0",x"78",x"c0",x"48"),
   263 => (x"4c",x"fd",x"87",x"c2"),
   264 => (x"fa",x"c3",x"4d",x"c1"),
   265 => (x"dd",x"de",x"ff",x"49"),
   266 => (x"c2",x"49",x"70",x"87"),
   267 => (x"d9",x"c0",x"02",x"99"),
   268 => (x"d9",x"ee",x"c2",x"87"),
   269 => (x"b7",x"c7",x"48",x"bf"),
   270 => (x"c9",x"c0",x"03",x"a8"),
   271 => (x"d9",x"ee",x"c2",x"87"),
   272 => (x"c0",x"78",x"c7",x"48"),
   273 => (x"4c",x"fc",x"87",x"c2"),
   274 => (x"b7",x"c0",x"4d",x"c1"),
   275 => (x"d3",x"c0",x"03",x"ac"),
   276 => (x"48",x"66",x"c4",x"87"),
   277 => (x"70",x"80",x"d8",x"c1"),
   278 => (x"02",x"bf",x"6e",x"7e"),
   279 => (x"4b",x"87",x"c5",x"c0"),
   280 => (x"0f",x"73",x"49",x"74"),
   281 => (x"f0",x"c3",x"1e",x"c0"),
   282 => (x"49",x"da",x"c1",x"1e"),
   283 => (x"c8",x"87",x"ca",x"f7"),
   284 => (x"02",x"98",x"70",x"86"),
   285 => (x"c2",x"87",x"d8",x"c0"),
   286 => (x"7e",x"bf",x"d9",x"ee"),
   287 => (x"91",x"cb",x"49",x"6e"),
   288 => (x"71",x"4a",x"66",x"c4"),
   289 => (x"c0",x"02",x"6a",x"82"),
   290 => (x"6e",x"4b",x"87",x"c5"),
   291 => (x"75",x"0f",x"73",x"49"),
   292 => (x"c8",x"c0",x"02",x"9d"),
   293 => (x"d9",x"ee",x"c2",x"87"),
   294 => (x"e0",x"f2",x"49",x"bf"),
   295 => (x"e4",x"d4",x"c2",x"87"),
   296 => (x"dd",x"c0",x"02",x"bf"),
   297 => (x"cb",x"c2",x"49",x"87"),
   298 => (x"02",x"98",x"70",x"87"),
   299 => (x"c2",x"87",x"d3",x"c0"),
   300 => (x"49",x"bf",x"d9",x"ee"),
   301 => (x"c0",x"87",x"c6",x"f2"),
   302 => (x"87",x"e6",x"f3",x"49"),
   303 => (x"48",x"e4",x"d4",x"c2"),
   304 => (x"8e",x"f8",x"78",x"c0"),
   305 => (x"0e",x"87",x"c0",x"f3"),
   306 => (x"5d",x"5c",x"5b",x"5e"),
   307 => (x"4c",x"71",x"1e",x"0e"),
   308 => (x"bf",x"d5",x"ee",x"c2"),
   309 => (x"a1",x"cd",x"c1",x"49"),
   310 => (x"81",x"d1",x"c1",x"4d"),
   311 => (x"9c",x"74",x"7e",x"69"),
   312 => (x"c4",x"87",x"cf",x"02"),
   313 => (x"7b",x"74",x"4b",x"a5"),
   314 => (x"bf",x"d5",x"ee",x"c2"),
   315 => (x"87",x"df",x"f2",x"49"),
   316 => (x"9c",x"74",x"7b",x"6e"),
   317 => (x"c0",x"87",x"c4",x"05"),
   318 => (x"c1",x"87",x"c2",x"4b"),
   319 => (x"f2",x"49",x"73",x"4b"),
   320 => (x"66",x"d4",x"87",x"e0"),
   321 => (x"49",x"87",x"c7",x"02"),
   322 => (x"4a",x"70",x"87",x"de"),
   323 => (x"4a",x"c0",x"87",x"c2"),
   324 => (x"5a",x"e8",x"d4",x"c2"),
   325 => (x"87",x"ef",x"f1",x"26"),
   326 => (x"00",x"00",x"00",x"00"),
   327 => (x"00",x"00",x"00",x"00"),
   328 => (x"00",x"00",x"00",x"00"),
   329 => (x"00",x"00",x"00",x"00"),
   330 => (x"ff",x"4a",x"71",x"1e"),
   331 => (x"72",x"49",x"bf",x"c8"),
   332 => (x"4f",x"26",x"48",x"a1"),
   333 => (x"bf",x"c8",x"ff",x"1e"),
   334 => (x"c0",x"c0",x"fe",x"89"),
   335 => (x"a9",x"c0",x"c0",x"c0"),
   336 => (x"c0",x"87",x"c4",x"01"),
   337 => (x"c1",x"87",x"c2",x"4a"),
   338 => (x"26",x"48",x"72",x"4a"),
   339 => (x"5b",x"5e",x"0e",x"4f"),
   340 => (x"71",x"0e",x"5d",x"5c"),
   341 => (x"4c",x"d4",x"ff",x"4b"),
   342 => (x"c0",x"48",x"66",x"d0"),
   343 => (x"ff",x"49",x"d6",x"78"),
   344 => (x"c3",x"87",x"db",x"db"),
   345 => (x"49",x"6c",x"7c",x"ff"),
   346 => (x"71",x"99",x"ff",x"c3"),
   347 => (x"f0",x"c3",x"49",x"4d"),
   348 => (x"a9",x"e0",x"c1",x"99"),
   349 => (x"c3",x"87",x"cb",x"05"),
   350 => (x"48",x"6c",x"7c",x"ff"),
   351 => (x"66",x"d0",x"98",x"c3"),
   352 => (x"ff",x"c3",x"78",x"08"),
   353 => (x"49",x"4a",x"6c",x"7c"),
   354 => (x"ff",x"c3",x"31",x"c8"),
   355 => (x"71",x"4a",x"6c",x"7c"),
   356 => (x"c8",x"49",x"72",x"b2"),
   357 => (x"7c",x"ff",x"c3",x"31"),
   358 => (x"b2",x"71",x"4a",x"6c"),
   359 => (x"31",x"c8",x"49",x"72"),
   360 => (x"6c",x"7c",x"ff",x"c3"),
   361 => (x"ff",x"b2",x"71",x"4a"),
   362 => (x"e0",x"c0",x"48",x"d0"),
   363 => (x"02",x"9b",x"73",x"78"),
   364 => (x"7b",x"72",x"87",x"c2"),
   365 => (x"4d",x"26",x"48",x"75"),
   366 => (x"4b",x"26",x"4c",x"26"),
   367 => (x"26",x"1e",x"4f",x"26"),
   368 => (x"5b",x"5e",x"0e",x"4f"),
   369 => (x"86",x"f8",x"0e",x"5c"),
   370 => (x"a6",x"c8",x"1e",x"76"),
   371 => (x"87",x"fd",x"fd",x"49"),
   372 => (x"4b",x"70",x"86",x"c4"),
   373 => (x"a8",x"c2",x"48",x"6e"),
   374 => (x"87",x"f0",x"c2",x"03"),
   375 => (x"f0",x"c3",x"4a",x"73"),
   376 => (x"aa",x"d0",x"c1",x"9a"),
   377 => (x"c1",x"87",x"c7",x"02"),
   378 => (x"c2",x"05",x"aa",x"e0"),
   379 => (x"49",x"73",x"87",x"de"),
   380 => (x"c3",x"02",x"99",x"c8"),
   381 => (x"87",x"c6",x"ff",x"87"),
   382 => (x"9c",x"c3",x"4c",x"73"),
   383 => (x"c1",x"05",x"ac",x"c2"),
   384 => (x"66",x"c4",x"87",x"c2"),
   385 => (x"71",x"31",x"c9",x"49"),
   386 => (x"4a",x"66",x"c4",x"1e"),
   387 => (x"ee",x"c2",x"92",x"d4"),
   388 => (x"81",x"72",x"49",x"dd"),
   389 => (x"87",x"fa",x"ce",x"fe"),
   390 => (x"d8",x"ff",x"49",x"d8"),
   391 => (x"c0",x"c8",x"87",x"e0"),
   392 => (x"fa",x"dc",x"c2",x"1e"),
   393 => (x"f5",x"ea",x"fd",x"49"),
   394 => (x"48",x"d0",x"ff",x"87"),
   395 => (x"c2",x"78",x"e0",x"c0"),
   396 => (x"cc",x"1e",x"fa",x"dc"),
   397 => (x"92",x"d4",x"4a",x"66"),
   398 => (x"49",x"dd",x"ee",x"c2"),
   399 => (x"cd",x"fe",x"81",x"72"),
   400 => (x"86",x"cc",x"87",x"c1"),
   401 => (x"c1",x"05",x"ac",x"c1"),
   402 => (x"66",x"c4",x"87",x"c2"),
   403 => (x"71",x"31",x"c9",x"49"),
   404 => (x"4a",x"66",x"c4",x"1e"),
   405 => (x"ee",x"c2",x"92",x"d4"),
   406 => (x"81",x"72",x"49",x"dd"),
   407 => (x"87",x"f2",x"cd",x"fe"),
   408 => (x"1e",x"fa",x"dc",x"c2"),
   409 => (x"d4",x"4a",x"66",x"c8"),
   410 => (x"dd",x"ee",x"c2",x"92"),
   411 => (x"fe",x"81",x"72",x"49"),
   412 => (x"d7",x"87",x"c1",x"cb"),
   413 => (x"c5",x"d7",x"ff",x"49"),
   414 => (x"1e",x"c0",x"c8",x"87"),
   415 => (x"49",x"fa",x"dc",x"c2"),
   416 => (x"87",x"f3",x"e8",x"fd"),
   417 => (x"d0",x"ff",x"86",x"cc"),
   418 => (x"78",x"e0",x"c0",x"48"),
   419 => (x"e7",x"fc",x"8e",x"f8"),
   420 => (x"5b",x"5e",x"0e",x"87"),
   421 => (x"1e",x"0e",x"5d",x"5c"),
   422 => (x"d4",x"ff",x"4d",x"71"),
   423 => (x"7e",x"66",x"d4",x"4c"),
   424 => (x"a8",x"b7",x"c3",x"48"),
   425 => (x"c0",x"87",x"c5",x"06"),
   426 => (x"87",x"e2",x"c1",x"48"),
   427 => (x"db",x"fe",x"49",x"75"),
   428 => (x"1e",x"75",x"87",x"ed"),
   429 => (x"d4",x"4b",x"66",x"c4"),
   430 => (x"dd",x"ee",x"c2",x"93"),
   431 => (x"fe",x"49",x"73",x"83"),
   432 => (x"c8",x"87",x"fd",x"c4"),
   433 => (x"ff",x"4b",x"6b",x"83"),
   434 => (x"e1",x"c8",x"48",x"d0"),
   435 => (x"73",x"7c",x"dd",x"78"),
   436 => (x"99",x"ff",x"c3",x"49"),
   437 => (x"49",x"73",x"7c",x"71"),
   438 => (x"c3",x"29",x"b7",x"c8"),
   439 => (x"7c",x"71",x"99",x"ff"),
   440 => (x"b7",x"d0",x"49",x"73"),
   441 => (x"99",x"ff",x"c3",x"29"),
   442 => (x"49",x"73",x"7c",x"71"),
   443 => (x"71",x"29",x"b7",x"d8"),
   444 => (x"7c",x"7c",x"c0",x"7c"),
   445 => (x"7c",x"7c",x"7c",x"7c"),
   446 => (x"7c",x"7c",x"7c",x"7c"),
   447 => (x"e0",x"c0",x"7c",x"7c"),
   448 => (x"1e",x"66",x"c4",x"78"),
   449 => (x"d5",x"ff",x"49",x"dc"),
   450 => (x"86",x"c8",x"87",x"d9"),
   451 => (x"fa",x"26",x"48",x"73"),
   452 => (x"fa",x"26",x"87",x"e4"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

