
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c8",x"ef",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c8",x"ef",x"c2"),
    14 => (x"48",x"d4",x"dc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e7",x"e3"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"49",x"72"),
    82 => (x"c2",x"7c",x"71",x"99"),
    83 => (x"05",x"bf",x"d4",x"dc"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"c3",x"29",x"d8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"d0",x"49",x"66",x"d0"),
    90 => (x"99",x"ff",x"c3",x"29"),
    91 => (x"66",x"d0",x"7c",x"71"),
    92 => (x"c3",x"29",x"c8",x"49"),
    93 => (x"7c",x"71",x"99",x"ff"),
    94 => (x"c3",x"49",x"66",x"d0"),
    95 => (x"7c",x"71",x"99",x"ff"),
    96 => (x"29",x"d0",x"49",x"72"),
    97 => (x"71",x"99",x"ff",x"c3"),
    98 => (x"c9",x"4b",x"6c",x"7c"),
    99 => (x"c3",x"4d",x"ff",x"f0"),
   100 => (x"d0",x"05",x"ab",x"ff"),
   101 => (x"7c",x"ff",x"c3",x"87"),
   102 => (x"8d",x"c1",x"4b",x"6c"),
   103 => (x"c3",x"87",x"c6",x"02"),
   104 => (x"f0",x"02",x"ab",x"ff"),
   105 => (x"fe",x"48",x"73",x"87"),
   106 => (x"c0",x"1e",x"87",x"c7"),
   107 => (x"48",x"d4",x"ff",x"49"),
   108 => (x"c1",x"78",x"ff",x"c3"),
   109 => (x"b7",x"c8",x"c3",x"81"),
   110 => (x"87",x"f1",x"04",x"a9"),
   111 => (x"73",x"1e",x"4f",x"26"),
   112 => (x"c4",x"87",x"e7",x"1e"),
   113 => (x"c0",x"4b",x"df",x"f8"),
   114 => (x"f0",x"ff",x"c0",x"1e"),
   115 => (x"fd",x"49",x"f7",x"c1"),
   116 => (x"86",x"c4",x"87",x"e7"),
   117 => (x"c0",x"05",x"a8",x"c1"),
   118 => (x"d4",x"ff",x"87",x"ea"),
   119 => (x"78",x"ff",x"c3",x"48"),
   120 => (x"c0",x"c0",x"c0",x"c1"),
   121 => (x"c0",x"1e",x"c0",x"c0"),
   122 => (x"e9",x"c1",x"f0",x"e1"),
   123 => (x"87",x"c9",x"fd",x"49"),
   124 => (x"98",x"70",x"86",x"c4"),
   125 => (x"ff",x"87",x"ca",x"05"),
   126 => (x"ff",x"c3",x"48",x"d4"),
   127 => (x"cb",x"48",x"c1",x"78"),
   128 => (x"87",x"e6",x"fe",x"87"),
   129 => (x"fe",x"05",x"8b",x"c1"),
   130 => (x"48",x"c0",x"87",x"fd"),
   131 => (x"1e",x"87",x"e6",x"fc"),
   132 => (x"d4",x"ff",x"1e",x"73"),
   133 => (x"78",x"ff",x"c3",x"48"),
   134 => (x"1e",x"c0",x"4b",x"d3"),
   135 => (x"c1",x"f0",x"ff",x"c0"),
   136 => (x"d4",x"fc",x"49",x"c1"),
   137 => (x"70",x"86",x"c4",x"87"),
   138 => (x"87",x"ca",x"05",x"98"),
   139 => (x"c3",x"48",x"d4",x"ff"),
   140 => (x"48",x"c1",x"78",x"ff"),
   141 => (x"f1",x"fd",x"87",x"cb"),
   142 => (x"05",x"8b",x"c1",x"87"),
   143 => (x"c0",x"87",x"db",x"ff"),
   144 => (x"87",x"f1",x"fb",x"48"),
   145 => (x"5c",x"5b",x"5e",x"0e"),
   146 => (x"4c",x"d4",x"ff",x"0e"),
   147 => (x"c6",x"87",x"db",x"fd"),
   148 => (x"e1",x"c0",x"1e",x"ea"),
   149 => (x"49",x"c8",x"c1",x"f0"),
   150 => (x"c4",x"87",x"de",x"fb"),
   151 => (x"02",x"a8",x"c1",x"86"),
   152 => (x"ea",x"fe",x"87",x"c8"),
   153 => (x"c1",x"48",x"c0",x"87"),
   154 => (x"da",x"fa",x"87",x"e2"),
   155 => (x"cf",x"49",x"70",x"87"),
   156 => (x"c6",x"99",x"ff",x"ff"),
   157 => (x"c8",x"02",x"a9",x"ea"),
   158 => (x"87",x"d3",x"fe",x"87"),
   159 => (x"cb",x"c1",x"48",x"c0"),
   160 => (x"7c",x"ff",x"c3",x"87"),
   161 => (x"fc",x"4b",x"f1",x"c0"),
   162 => (x"98",x"70",x"87",x"f4"),
   163 => (x"87",x"eb",x"c0",x"02"),
   164 => (x"ff",x"c0",x"1e",x"c0"),
   165 => (x"49",x"fa",x"c1",x"f0"),
   166 => (x"c4",x"87",x"de",x"fa"),
   167 => (x"05",x"98",x"70",x"86"),
   168 => (x"ff",x"c3",x"87",x"d9"),
   169 => (x"c3",x"49",x"6c",x"7c"),
   170 => (x"7c",x"7c",x"7c",x"ff"),
   171 => (x"99",x"c0",x"c1",x"7c"),
   172 => (x"c1",x"87",x"c4",x"02"),
   173 => (x"c0",x"87",x"d5",x"48"),
   174 => (x"c2",x"87",x"d1",x"48"),
   175 => (x"87",x"c4",x"05",x"ab"),
   176 => (x"87",x"c8",x"48",x"c0"),
   177 => (x"fe",x"05",x"8b",x"c1"),
   178 => (x"48",x"c0",x"87",x"fd"),
   179 => (x"1e",x"87",x"e4",x"f9"),
   180 => (x"dc",x"c2",x"1e",x"73"),
   181 => (x"78",x"c1",x"48",x"d4"),
   182 => (x"d0",x"ff",x"4b",x"c7"),
   183 => (x"fb",x"78",x"c2",x"48"),
   184 => (x"d0",x"ff",x"87",x"c8"),
   185 => (x"c0",x"78",x"c3",x"48"),
   186 => (x"d0",x"e5",x"c0",x"1e"),
   187 => (x"f9",x"49",x"c0",x"c1"),
   188 => (x"86",x"c4",x"87",x"c7"),
   189 => (x"c1",x"05",x"a8",x"c1"),
   190 => (x"ab",x"c2",x"4b",x"87"),
   191 => (x"c0",x"87",x"c5",x"05"),
   192 => (x"87",x"f9",x"c0",x"48"),
   193 => (x"ff",x"05",x"8b",x"c1"),
   194 => (x"f7",x"fc",x"87",x"d0"),
   195 => (x"d8",x"dc",x"c2",x"87"),
   196 => (x"05",x"98",x"70",x"58"),
   197 => (x"1e",x"c1",x"87",x"cd"),
   198 => (x"c1",x"f0",x"ff",x"c0"),
   199 => (x"d8",x"f8",x"49",x"d0"),
   200 => (x"ff",x"86",x"c4",x"87"),
   201 => (x"ff",x"c3",x"48",x"d4"),
   202 => (x"87",x"de",x"c4",x"78"),
   203 => (x"58",x"dc",x"dc",x"c2"),
   204 => (x"c2",x"48",x"d0",x"ff"),
   205 => (x"48",x"d4",x"ff",x"78"),
   206 => (x"c1",x"78",x"ff",x"c3"),
   207 => (x"87",x"f5",x"f7",x"48"),
   208 => (x"5c",x"5b",x"5e",x"0e"),
   209 => (x"4a",x"71",x"0e",x"5d"),
   210 => (x"ff",x"4d",x"ff",x"c3"),
   211 => (x"7c",x"75",x"4c",x"d4"),
   212 => (x"c4",x"48",x"d0",x"ff"),
   213 => (x"7c",x"75",x"78",x"c3"),
   214 => (x"ff",x"c0",x"1e",x"72"),
   215 => (x"49",x"d8",x"c1",x"f0"),
   216 => (x"c4",x"87",x"d6",x"f7"),
   217 => (x"02",x"98",x"70",x"86"),
   218 => (x"48",x"c1",x"87",x"c5"),
   219 => (x"75",x"87",x"f0",x"c0"),
   220 => (x"7c",x"fe",x"c3",x"7c"),
   221 => (x"d4",x"1e",x"c0",x"c8"),
   222 => (x"fa",x"f4",x"49",x"66"),
   223 => (x"75",x"86",x"c4",x"87"),
   224 => (x"75",x"7c",x"75",x"7c"),
   225 => (x"e0",x"da",x"d8",x"7c"),
   226 => (x"6c",x"7c",x"75",x"4b"),
   227 => (x"c5",x"05",x"99",x"49"),
   228 => (x"05",x"8b",x"c1",x"87"),
   229 => (x"7c",x"75",x"87",x"f3"),
   230 => (x"c2",x"48",x"d0",x"ff"),
   231 => (x"f6",x"48",x"c0",x"78"),
   232 => (x"5e",x"0e",x"87",x"cf"),
   233 => (x"0e",x"5d",x"5c",x"5b"),
   234 => (x"4c",x"c0",x"4b",x"71"),
   235 => (x"df",x"cd",x"ee",x"c5"),
   236 => (x"48",x"d4",x"ff",x"4a"),
   237 => (x"68",x"78",x"ff",x"c3"),
   238 => (x"a9",x"fe",x"c3",x"49"),
   239 => (x"87",x"fd",x"c0",x"05"),
   240 => (x"9b",x"73",x"4d",x"70"),
   241 => (x"d0",x"87",x"cc",x"02"),
   242 => (x"49",x"73",x"1e",x"66"),
   243 => (x"c4",x"87",x"cf",x"f4"),
   244 => (x"ff",x"87",x"d6",x"86"),
   245 => (x"d1",x"c4",x"48",x"d0"),
   246 => (x"7d",x"ff",x"c3",x"78"),
   247 => (x"c1",x"48",x"66",x"d0"),
   248 => (x"58",x"a6",x"d4",x"88"),
   249 => (x"f0",x"05",x"98",x"70"),
   250 => (x"48",x"d4",x"ff",x"87"),
   251 => (x"78",x"78",x"ff",x"c3"),
   252 => (x"c5",x"05",x"9b",x"73"),
   253 => (x"48",x"d0",x"ff",x"87"),
   254 => (x"4a",x"c1",x"78",x"d0"),
   255 => (x"05",x"8a",x"c1",x"4c"),
   256 => (x"74",x"87",x"ee",x"fe"),
   257 => (x"87",x"e9",x"f4",x"48"),
   258 => (x"71",x"1e",x"73",x"1e"),
   259 => (x"ff",x"4b",x"c0",x"4a"),
   260 => (x"ff",x"c3",x"48",x"d4"),
   261 => (x"48",x"d0",x"ff",x"78"),
   262 => (x"ff",x"78",x"c3",x"c4"),
   263 => (x"ff",x"c3",x"48",x"d4"),
   264 => (x"c0",x"1e",x"72",x"78"),
   265 => (x"d1",x"c1",x"f0",x"ff"),
   266 => (x"87",x"cd",x"f4",x"49"),
   267 => (x"98",x"70",x"86",x"c4"),
   268 => (x"c8",x"87",x"d2",x"05"),
   269 => (x"66",x"cc",x"1e",x"c0"),
   270 => (x"87",x"e6",x"fd",x"49"),
   271 => (x"4b",x"70",x"86",x"c4"),
   272 => (x"c2",x"48",x"d0",x"ff"),
   273 => (x"f3",x"48",x"73",x"78"),
   274 => (x"5e",x"0e",x"87",x"eb"),
   275 => (x"0e",x"5d",x"5c",x"5b"),
   276 => (x"ff",x"c0",x"1e",x"c0"),
   277 => (x"49",x"c9",x"c1",x"f0"),
   278 => (x"d2",x"87",x"de",x"f3"),
   279 => (x"dc",x"dc",x"c2",x"1e"),
   280 => (x"87",x"fe",x"fc",x"49"),
   281 => (x"4c",x"c0",x"86",x"c8"),
   282 => (x"b7",x"d2",x"84",x"c1"),
   283 => (x"87",x"f8",x"04",x"ac"),
   284 => (x"97",x"dc",x"dc",x"c2"),
   285 => (x"c0",x"c3",x"49",x"bf"),
   286 => (x"a9",x"c0",x"c1",x"99"),
   287 => (x"87",x"e7",x"c0",x"05"),
   288 => (x"97",x"e3",x"dc",x"c2"),
   289 => (x"31",x"d0",x"49",x"bf"),
   290 => (x"97",x"e4",x"dc",x"c2"),
   291 => (x"32",x"c8",x"4a",x"bf"),
   292 => (x"dc",x"c2",x"b1",x"72"),
   293 => (x"4a",x"bf",x"97",x"e5"),
   294 => (x"cf",x"4c",x"71",x"b1"),
   295 => (x"9c",x"ff",x"ff",x"ff"),
   296 => (x"34",x"ca",x"84",x"c1"),
   297 => (x"c2",x"87",x"e7",x"c1"),
   298 => (x"bf",x"97",x"e5",x"dc"),
   299 => (x"c6",x"31",x"c1",x"49"),
   300 => (x"e6",x"dc",x"c2",x"99"),
   301 => (x"c7",x"4a",x"bf",x"97"),
   302 => (x"b1",x"72",x"2a",x"b7"),
   303 => (x"97",x"e1",x"dc",x"c2"),
   304 => (x"cf",x"4d",x"4a",x"bf"),
   305 => (x"e2",x"dc",x"c2",x"9d"),
   306 => (x"c3",x"4a",x"bf",x"97"),
   307 => (x"c2",x"32",x"ca",x"9a"),
   308 => (x"bf",x"97",x"e3",x"dc"),
   309 => (x"73",x"33",x"c2",x"4b"),
   310 => (x"e4",x"dc",x"c2",x"b2"),
   311 => (x"c3",x"4b",x"bf",x"97"),
   312 => (x"b7",x"c6",x"9b",x"c0"),
   313 => (x"c2",x"b2",x"73",x"2b"),
   314 => (x"71",x"48",x"c1",x"81"),
   315 => (x"c1",x"49",x"70",x"30"),
   316 => (x"70",x"30",x"75",x"48"),
   317 => (x"c1",x"4c",x"72",x"4d"),
   318 => (x"c8",x"94",x"71",x"84"),
   319 => (x"06",x"ad",x"b7",x"c0"),
   320 => (x"34",x"c1",x"87",x"cc"),
   321 => (x"c0",x"c8",x"2d",x"b7"),
   322 => (x"ff",x"01",x"ad",x"b7"),
   323 => (x"48",x"74",x"87",x"f4"),
   324 => (x"0e",x"87",x"de",x"f0"),
   325 => (x"5d",x"5c",x"5b",x"5e"),
   326 => (x"c2",x"86",x"f8",x"0e"),
   327 => (x"c0",x"48",x"c2",x"e5"),
   328 => (x"fa",x"dc",x"c2",x"78"),
   329 => (x"fb",x"49",x"c0",x"1e"),
   330 => (x"86",x"c4",x"87",x"de"),
   331 => (x"c5",x"05",x"98",x"70"),
   332 => (x"c9",x"48",x"c0",x"87"),
   333 => (x"4d",x"c0",x"87",x"ce"),
   334 => (x"f2",x"c0",x"7e",x"c1"),
   335 => (x"c2",x"49",x"bf",x"ed"),
   336 => (x"71",x"4a",x"f0",x"dd"),
   337 => (x"e0",x"ec",x"4b",x"c8"),
   338 => (x"05",x"98",x"70",x"87"),
   339 => (x"7e",x"c0",x"87",x"c2"),
   340 => (x"bf",x"e9",x"f2",x"c0"),
   341 => (x"cc",x"de",x"c2",x"49"),
   342 => (x"4b",x"c8",x"71",x"4a"),
   343 => (x"70",x"87",x"ca",x"ec"),
   344 => (x"87",x"c2",x"05",x"98"),
   345 => (x"02",x"6e",x"7e",x"c0"),
   346 => (x"c2",x"87",x"fd",x"c0"),
   347 => (x"4d",x"bf",x"c0",x"e4"),
   348 => (x"9f",x"f8",x"e4",x"c2"),
   349 => (x"c5",x"48",x"7e",x"bf"),
   350 => (x"05",x"a8",x"ea",x"d6"),
   351 => (x"e4",x"c2",x"87",x"c7"),
   352 => (x"ce",x"4d",x"bf",x"c0"),
   353 => (x"ca",x"48",x"6e",x"87"),
   354 => (x"02",x"a8",x"d5",x"e9"),
   355 => (x"48",x"c0",x"87",x"c5"),
   356 => (x"c2",x"87",x"f1",x"c7"),
   357 => (x"75",x"1e",x"fa",x"dc"),
   358 => (x"87",x"ec",x"f9",x"49"),
   359 => (x"98",x"70",x"86",x"c4"),
   360 => (x"c0",x"87",x"c5",x"05"),
   361 => (x"87",x"dc",x"c7",x"48"),
   362 => (x"bf",x"e9",x"f2",x"c0"),
   363 => (x"cc",x"de",x"c2",x"49"),
   364 => (x"4b",x"c8",x"71",x"4a"),
   365 => (x"70",x"87",x"f2",x"ea"),
   366 => (x"87",x"c8",x"05",x"98"),
   367 => (x"48",x"c2",x"e5",x"c2"),
   368 => (x"87",x"da",x"78",x"c1"),
   369 => (x"bf",x"ed",x"f2",x"c0"),
   370 => (x"f0",x"dd",x"c2",x"49"),
   371 => (x"4b",x"c8",x"71",x"4a"),
   372 => (x"70",x"87",x"d6",x"ea"),
   373 => (x"c5",x"c0",x"02",x"98"),
   374 => (x"c6",x"48",x"c0",x"87"),
   375 => (x"e4",x"c2",x"87",x"e6"),
   376 => (x"49",x"bf",x"97",x"f8"),
   377 => (x"05",x"a9",x"d5",x"c1"),
   378 => (x"c2",x"87",x"cd",x"c0"),
   379 => (x"bf",x"97",x"f9",x"e4"),
   380 => (x"a9",x"ea",x"c2",x"49"),
   381 => (x"87",x"c5",x"c0",x"02"),
   382 => (x"c7",x"c6",x"48",x"c0"),
   383 => (x"fa",x"dc",x"c2",x"87"),
   384 => (x"48",x"7e",x"bf",x"97"),
   385 => (x"02",x"a8",x"e9",x"c3"),
   386 => (x"6e",x"87",x"ce",x"c0"),
   387 => (x"a8",x"eb",x"c3",x"48"),
   388 => (x"87",x"c5",x"c0",x"02"),
   389 => (x"eb",x"c5",x"48",x"c0"),
   390 => (x"c5",x"dd",x"c2",x"87"),
   391 => (x"99",x"49",x"bf",x"97"),
   392 => (x"87",x"cc",x"c0",x"05"),
   393 => (x"97",x"c6",x"dd",x"c2"),
   394 => (x"a9",x"c2",x"49",x"bf"),
   395 => (x"87",x"c5",x"c0",x"02"),
   396 => (x"cf",x"c5",x"48",x"c0"),
   397 => (x"c7",x"dd",x"c2",x"87"),
   398 => (x"c2",x"48",x"bf",x"97"),
   399 => (x"70",x"58",x"fe",x"e4"),
   400 => (x"88",x"c1",x"48",x"4c"),
   401 => (x"58",x"c2",x"e5",x"c2"),
   402 => (x"97",x"c8",x"dd",x"c2"),
   403 => (x"81",x"75",x"49",x"bf"),
   404 => (x"97",x"c9",x"dd",x"c2"),
   405 => (x"32",x"c8",x"4a",x"bf"),
   406 => (x"c2",x"7e",x"a1",x"72"),
   407 => (x"6e",x"48",x"cf",x"e9"),
   408 => (x"ca",x"dd",x"c2",x"78"),
   409 => (x"c8",x"48",x"bf",x"97"),
   410 => (x"e5",x"c2",x"58",x"a6"),
   411 => (x"c2",x"02",x"bf",x"c2"),
   412 => (x"f2",x"c0",x"87",x"d4"),
   413 => (x"c2",x"49",x"bf",x"e9"),
   414 => (x"71",x"4a",x"cc",x"de"),
   415 => (x"e8",x"e7",x"4b",x"c8"),
   416 => (x"02",x"98",x"70",x"87"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"f8",x"c3",x"48"),
   419 => (x"bf",x"fa",x"e4",x"c2"),
   420 => (x"e3",x"e9",x"c2",x"4c"),
   421 => (x"df",x"dd",x"c2",x"5c"),
   422 => (x"c8",x"49",x"bf",x"97"),
   423 => (x"de",x"dd",x"c2",x"31"),
   424 => (x"a1",x"4a",x"bf",x"97"),
   425 => (x"e0",x"dd",x"c2",x"49"),
   426 => (x"d0",x"4a",x"bf",x"97"),
   427 => (x"49",x"a1",x"72",x"32"),
   428 => (x"97",x"e1",x"dd",x"c2"),
   429 => (x"32",x"d8",x"4a",x"bf"),
   430 => (x"c4",x"49",x"a1",x"72"),
   431 => (x"e9",x"c2",x"91",x"66"),
   432 => (x"c2",x"81",x"bf",x"cf"),
   433 => (x"c2",x"59",x"d7",x"e9"),
   434 => (x"bf",x"97",x"e7",x"dd"),
   435 => (x"c2",x"32",x"c8",x"4a"),
   436 => (x"bf",x"97",x"e6",x"dd"),
   437 => (x"c2",x"4a",x"a2",x"4b"),
   438 => (x"bf",x"97",x"e8",x"dd"),
   439 => (x"73",x"33",x"d0",x"4b"),
   440 => (x"dd",x"c2",x"4a",x"a2"),
   441 => (x"4b",x"bf",x"97",x"e9"),
   442 => (x"33",x"d8",x"9b",x"cf"),
   443 => (x"c2",x"4a",x"a2",x"73"),
   444 => (x"c2",x"5a",x"db",x"e9"),
   445 => (x"4a",x"bf",x"d7",x"e9"),
   446 => (x"92",x"74",x"8a",x"c2"),
   447 => (x"48",x"db",x"e9",x"c2"),
   448 => (x"c1",x"78",x"a1",x"72"),
   449 => (x"dd",x"c2",x"87",x"ca"),
   450 => (x"49",x"bf",x"97",x"cc"),
   451 => (x"dd",x"c2",x"31",x"c8"),
   452 => (x"4a",x"bf",x"97",x"cb"),
   453 => (x"e5",x"c2",x"49",x"a1"),
   454 => (x"e5",x"c2",x"59",x"ca"),
   455 => (x"c5",x"49",x"bf",x"c6"),
   456 => (x"81",x"ff",x"c7",x"31"),
   457 => (x"e9",x"c2",x"29",x"c9"),
   458 => (x"dd",x"c2",x"59",x"e3"),
   459 => (x"4a",x"bf",x"97",x"d1"),
   460 => (x"dd",x"c2",x"32",x"c8"),
   461 => (x"4b",x"bf",x"97",x"d0"),
   462 => (x"66",x"c4",x"4a",x"a2"),
   463 => (x"c2",x"82",x"6e",x"92"),
   464 => (x"c2",x"5a",x"df",x"e9"),
   465 => (x"c0",x"48",x"d7",x"e9"),
   466 => (x"d3",x"e9",x"c2",x"78"),
   467 => (x"78",x"a1",x"72",x"48"),
   468 => (x"48",x"e3",x"e9",x"c2"),
   469 => (x"bf",x"d7",x"e9",x"c2"),
   470 => (x"e7",x"e9",x"c2",x"78"),
   471 => (x"db",x"e9",x"c2",x"48"),
   472 => (x"e5",x"c2",x"78",x"bf"),
   473 => (x"c0",x"02",x"bf",x"c2"),
   474 => (x"48",x"74",x"87",x"c9"),
   475 => (x"7e",x"70",x"30",x"c4"),
   476 => (x"c2",x"87",x"c9",x"c0"),
   477 => (x"48",x"bf",x"df",x"e9"),
   478 => (x"7e",x"70",x"30",x"c4"),
   479 => (x"48",x"c6",x"e5",x"c2"),
   480 => (x"48",x"c1",x"78",x"6e"),
   481 => (x"4d",x"26",x"8e",x"f8"),
   482 => (x"4b",x"26",x"4c",x"26"),
   483 => (x"5e",x"0e",x"4f",x"26"),
   484 => (x"0e",x"5d",x"5c",x"5b"),
   485 => (x"e5",x"c2",x"4a",x"71"),
   486 => (x"cb",x"02",x"bf",x"c2"),
   487 => (x"c7",x"4b",x"72",x"87"),
   488 => (x"c1",x"4c",x"72",x"2b"),
   489 => (x"87",x"c9",x"9c",x"ff"),
   490 => (x"2b",x"c8",x"4b",x"72"),
   491 => (x"ff",x"c3",x"4c",x"72"),
   492 => (x"cf",x"e9",x"c2",x"9c"),
   493 => (x"f2",x"c0",x"83",x"bf"),
   494 => (x"02",x"ab",x"bf",x"e5"),
   495 => (x"f2",x"c0",x"87",x"d9"),
   496 => (x"dc",x"c2",x"5b",x"e9"),
   497 => (x"49",x"73",x"1e",x"fa"),
   498 => (x"c4",x"87",x"fd",x"f0"),
   499 => (x"05",x"98",x"70",x"86"),
   500 => (x"48",x"c0",x"87",x"c5"),
   501 => (x"c2",x"87",x"e6",x"c0"),
   502 => (x"02",x"bf",x"c2",x"e5"),
   503 => (x"49",x"74",x"87",x"d2"),
   504 => (x"dc",x"c2",x"91",x"c4"),
   505 => (x"4d",x"69",x"81",x"fa"),
   506 => (x"ff",x"ff",x"ff",x"cf"),
   507 => (x"87",x"cb",x"9d",x"ff"),
   508 => (x"91",x"c2",x"49",x"74"),
   509 => (x"81",x"fa",x"dc",x"c2"),
   510 => (x"75",x"4d",x"69",x"9f"),
   511 => (x"87",x"c6",x"fe",x"48"),
   512 => (x"5c",x"5b",x"5e",x"0e"),
   513 => (x"86",x"f8",x"0e",x"5d"),
   514 => (x"05",x"9c",x"4c",x"71"),
   515 => (x"48",x"c0",x"87",x"c5"),
   516 => (x"c8",x"87",x"c2",x"c3"),
   517 => (x"48",x"6e",x"7e",x"a4"),
   518 => (x"66",x"d8",x"78",x"c0"),
   519 => (x"d8",x"87",x"c7",x"02"),
   520 => (x"05",x"bf",x"97",x"66"),
   521 => (x"48",x"c0",x"87",x"c5"),
   522 => (x"c0",x"87",x"ea",x"c2"),
   523 => (x"49",x"49",x"c1",x"1e"),
   524 => (x"c4",x"87",x"d7",x"ca"),
   525 => (x"9d",x"4d",x"70",x"86"),
   526 => (x"87",x"c2",x"c1",x"02"),
   527 => (x"4a",x"ca",x"e5",x"c2"),
   528 => (x"e0",x"49",x"66",x"d8"),
   529 => (x"98",x"70",x"87",x"c8"),
   530 => (x"87",x"f2",x"c0",x"02"),
   531 => (x"66",x"d8",x"4a",x"75"),
   532 => (x"e0",x"4b",x"cb",x"49"),
   533 => (x"98",x"70",x"87",x"ed"),
   534 => (x"87",x"e2",x"c0",x"02"),
   535 => (x"9d",x"75",x"1e",x"c0"),
   536 => (x"c8",x"87",x"c7",x"02"),
   537 => (x"78",x"c0",x"48",x"a6"),
   538 => (x"a6",x"c8",x"87",x"c5"),
   539 => (x"c8",x"78",x"c1",x"48"),
   540 => (x"d5",x"c9",x"49",x"66"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"fe",x"05",x"9d",x"4d"),
   543 => (x"9d",x"75",x"87",x"fe"),
   544 => (x"87",x"cf",x"c1",x"02"),
   545 => (x"6e",x"49",x"a5",x"dc"),
   546 => (x"da",x"78",x"69",x"48"),
   547 => (x"a6",x"c4",x"49",x"a5"),
   548 => (x"78",x"a4",x"c4",x"48"),
   549 => (x"c4",x"48",x"69",x"9f"),
   550 => (x"c2",x"78",x"08",x"66"),
   551 => (x"02",x"bf",x"c2",x"e5"),
   552 => (x"a5",x"d4",x"87",x"d2"),
   553 => (x"49",x"69",x"9f",x"49"),
   554 => (x"99",x"ff",x"ff",x"c0"),
   555 => (x"30",x"d0",x"48",x"71"),
   556 => (x"87",x"c2",x"7e",x"70"),
   557 => (x"49",x"6e",x"7e",x"c0"),
   558 => (x"bf",x"66",x"c4",x"48"),
   559 => (x"08",x"66",x"c4",x"80"),
   560 => (x"cc",x"7c",x"c0",x"78"),
   561 => (x"66",x"c4",x"49",x"a4"),
   562 => (x"a4",x"d0",x"79",x"bf"),
   563 => (x"c1",x"79",x"c0",x"49"),
   564 => (x"c0",x"87",x"c2",x"48"),
   565 => (x"fa",x"8e",x"f8",x"48"),
   566 => (x"5e",x"0e",x"87",x"ec"),
   567 => (x"0e",x"5d",x"5c",x"5b"),
   568 => (x"02",x"9c",x"4c",x"71"),
   569 => (x"c8",x"87",x"ca",x"c1"),
   570 => (x"02",x"69",x"49",x"a4"),
   571 => (x"d0",x"87",x"c2",x"c1"),
   572 => (x"49",x"6c",x"4a",x"66"),
   573 => (x"5a",x"a6",x"d4",x"82"),
   574 => (x"b9",x"4d",x"66",x"d0"),
   575 => (x"bf",x"fe",x"e4",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"02",x"99",x"71",x"99"),
   578 => (x"c4",x"87",x"e4",x"c0"),
   579 => (x"49",x"6b",x"4b",x"a4"),
   580 => (x"70",x"87",x"fb",x"f9"),
   581 => (x"fa",x"e4",x"c2",x"7b"),
   582 => (x"81",x"6c",x"49",x"bf"),
   583 => (x"b9",x"75",x"7c",x"71"),
   584 => (x"bf",x"fe",x"e4",x"c2"),
   585 => (x"72",x"ba",x"ff",x"4a"),
   586 => (x"05",x"99",x"71",x"99"),
   587 => (x"75",x"87",x"dc",x"ff"),
   588 => (x"87",x"d2",x"f9",x"7c"),
   589 => (x"71",x"1e",x"73",x"1e"),
   590 => (x"c7",x"02",x"9b",x"4b"),
   591 => (x"49",x"a3",x"c8",x"87"),
   592 => (x"87",x"c5",x"05",x"69"),
   593 => (x"f7",x"c0",x"48",x"c0"),
   594 => (x"d3",x"e9",x"c2",x"87"),
   595 => (x"a3",x"c4",x"4a",x"bf"),
   596 => (x"c2",x"49",x"69",x"49"),
   597 => (x"fa",x"e4",x"c2",x"89"),
   598 => (x"a2",x"71",x"91",x"bf"),
   599 => (x"fe",x"e4",x"c2",x"4a"),
   600 => (x"99",x"6b",x"49",x"bf"),
   601 => (x"c0",x"4a",x"a2",x"71"),
   602 => (x"c8",x"5a",x"e9",x"f2"),
   603 => (x"49",x"72",x"1e",x"66"),
   604 => (x"c4",x"87",x"d5",x"ea"),
   605 => (x"05",x"98",x"70",x"86"),
   606 => (x"48",x"c0",x"87",x"c4"),
   607 => (x"48",x"c1",x"87",x"c2"),
   608 => (x"1e",x"87",x"c7",x"f8"),
   609 => (x"4b",x"71",x"1e",x"73"),
   610 => (x"87",x"c7",x"02",x"9b"),
   611 => (x"69",x"49",x"a3",x"c8"),
   612 => (x"c0",x"87",x"c5",x"05"),
   613 => (x"87",x"f7",x"c0",x"48"),
   614 => (x"bf",x"d3",x"e9",x"c2"),
   615 => (x"49",x"a3",x"c4",x"4a"),
   616 => (x"89",x"c2",x"49",x"69"),
   617 => (x"bf",x"fa",x"e4",x"c2"),
   618 => (x"4a",x"a2",x"71",x"91"),
   619 => (x"bf",x"fe",x"e4",x"c2"),
   620 => (x"71",x"99",x"6b",x"49"),
   621 => (x"f2",x"c0",x"4a",x"a2"),
   622 => (x"66",x"c8",x"5a",x"e9"),
   623 => (x"e5",x"49",x"72",x"1e"),
   624 => (x"86",x"c4",x"87",x"fe"),
   625 => (x"c4",x"05",x"98",x"70"),
   626 => (x"c2",x"48",x"c0",x"87"),
   627 => (x"f6",x"48",x"c1",x"87"),
   628 => (x"5e",x"0e",x"87",x"f8"),
   629 => (x"0e",x"5d",x"5c",x"5b"),
   630 => (x"d4",x"4b",x"71",x"1e"),
   631 => (x"9b",x"73",x"4d",x"66"),
   632 => (x"87",x"cc",x"c1",x"02"),
   633 => (x"69",x"49",x"a3",x"c8"),
   634 => (x"87",x"c4",x"c1",x"02"),
   635 => (x"c2",x"4c",x"a3",x"d0"),
   636 => (x"49",x"bf",x"fe",x"e4"),
   637 => (x"4a",x"6c",x"b9",x"ff"),
   638 => (x"66",x"d4",x"7e",x"99"),
   639 => (x"87",x"cd",x"06",x"a9"),
   640 => (x"cc",x"7c",x"7b",x"c0"),
   641 => (x"a3",x"c4",x"4a",x"a3"),
   642 => (x"ca",x"79",x"6a",x"49"),
   643 => (x"f8",x"49",x"72",x"87"),
   644 => (x"66",x"d4",x"99",x"c0"),
   645 => (x"75",x"8d",x"71",x"4d"),
   646 => (x"71",x"29",x"c9",x"49"),
   647 => (x"fa",x"49",x"73",x"1e"),
   648 => (x"dc",x"c2",x"87",x"f8"),
   649 => (x"49",x"73",x"1e",x"fa"),
   650 => (x"c8",x"87",x"c9",x"fc"),
   651 => (x"7c",x"66",x"d4",x"86"),
   652 => (x"87",x"d2",x"f5",x"26"),
   653 => (x"71",x"1e",x"73",x"1e"),
   654 => (x"c0",x"02",x"9b",x"4b"),
   655 => (x"e9",x"c2",x"87",x"e4"),
   656 => (x"4a",x"73",x"5b",x"e7"),
   657 => (x"e4",x"c2",x"8a",x"c2"),
   658 => (x"92",x"49",x"bf",x"fa"),
   659 => (x"bf",x"d3",x"e9",x"c2"),
   660 => (x"c2",x"80",x"72",x"48"),
   661 => (x"71",x"58",x"eb",x"e9"),
   662 => (x"c2",x"30",x"c4",x"48"),
   663 => (x"c0",x"58",x"ca",x"e5"),
   664 => (x"e9",x"c2",x"87",x"ed"),
   665 => (x"e9",x"c2",x"48",x"e3"),
   666 => (x"c2",x"78",x"bf",x"d7"),
   667 => (x"c2",x"48",x"e7",x"e9"),
   668 => (x"78",x"bf",x"db",x"e9"),
   669 => (x"bf",x"c2",x"e5",x"c2"),
   670 => (x"c2",x"87",x"c9",x"02"),
   671 => (x"49",x"bf",x"fa",x"e4"),
   672 => (x"87",x"c7",x"31",x"c4"),
   673 => (x"bf",x"df",x"e9",x"c2"),
   674 => (x"c2",x"31",x"c4",x"49"),
   675 => (x"f3",x"59",x"ca",x"e5"),
   676 => (x"5e",x"0e",x"87",x"f8"),
   677 => (x"71",x"0e",x"5c",x"5b"),
   678 => (x"72",x"4b",x"c0",x"4a"),
   679 => (x"e1",x"c0",x"02",x"9a"),
   680 => (x"49",x"a2",x"da",x"87"),
   681 => (x"c2",x"4b",x"69",x"9f"),
   682 => (x"02",x"bf",x"c2",x"e5"),
   683 => (x"a2",x"d4",x"87",x"cf"),
   684 => (x"49",x"69",x"9f",x"49"),
   685 => (x"ff",x"ff",x"c0",x"4c"),
   686 => (x"c2",x"34",x"d0",x"9c"),
   687 => (x"74",x"4c",x"c0",x"87"),
   688 => (x"49",x"73",x"b3",x"49"),
   689 => (x"f2",x"87",x"ed",x"fd"),
   690 => (x"5e",x"0e",x"87",x"fe"),
   691 => (x"0e",x"5d",x"5c",x"5b"),
   692 => (x"4a",x"71",x"86",x"f4"),
   693 => (x"9a",x"72",x"7e",x"c0"),
   694 => (x"c2",x"87",x"d8",x"02"),
   695 => (x"c0",x"48",x"f6",x"dc"),
   696 => (x"ee",x"dc",x"c2",x"78"),
   697 => (x"e7",x"e9",x"c2",x"48"),
   698 => (x"dc",x"c2",x"78",x"bf"),
   699 => (x"e9",x"c2",x"48",x"f2"),
   700 => (x"c2",x"78",x"bf",x"e3"),
   701 => (x"c0",x"48",x"d7",x"e5"),
   702 => (x"c6",x"e5",x"c2",x"50"),
   703 => (x"dc",x"c2",x"49",x"bf"),
   704 => (x"71",x"4a",x"bf",x"f6"),
   705 => (x"c9",x"c4",x"03",x"aa"),
   706 => (x"cf",x"49",x"72",x"87"),
   707 => (x"e9",x"c0",x"05",x"99"),
   708 => (x"e5",x"f2",x"c0",x"87"),
   709 => (x"ee",x"dc",x"c2",x"48"),
   710 => (x"dc",x"c2",x"78",x"bf"),
   711 => (x"dc",x"c2",x"1e",x"fa"),
   712 => (x"c2",x"49",x"bf",x"ee"),
   713 => (x"c1",x"48",x"ee",x"dc"),
   714 => (x"e3",x"71",x"78",x"a1"),
   715 => (x"86",x"c4",x"87",x"da"),
   716 => (x"48",x"e1",x"f2",x"c0"),
   717 => (x"78",x"fa",x"dc",x"c2"),
   718 => (x"f2",x"c0",x"87",x"cc"),
   719 => (x"c0",x"48",x"bf",x"e1"),
   720 => (x"f2",x"c0",x"80",x"e0"),
   721 => (x"dc",x"c2",x"58",x"e5"),
   722 => (x"c1",x"48",x"bf",x"f6"),
   723 => (x"fa",x"dc",x"c2",x"80"),
   724 => (x"0c",x"a1",x"27",x"58"),
   725 => (x"97",x"bf",x"00",x"00"),
   726 => (x"02",x"9d",x"4d",x"bf"),
   727 => (x"c3",x"87",x"e3",x"c2"),
   728 => (x"c2",x"02",x"ad",x"e5"),
   729 => (x"f2",x"c0",x"87",x"dc"),
   730 => (x"cb",x"4b",x"bf",x"e1"),
   731 => (x"4c",x"11",x"49",x"a3"),
   732 => (x"c1",x"05",x"ac",x"cf"),
   733 => (x"49",x"75",x"87",x"d2"),
   734 => (x"89",x"c1",x"99",x"df"),
   735 => (x"e5",x"c2",x"91",x"cd"),
   736 => (x"a3",x"c1",x"81",x"ca"),
   737 => (x"c3",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"c5"),
   740 => (x"4a",x"a3",x"c7",x"51"),
   741 => (x"a3",x"c9",x"51",x"12"),
   742 => (x"ce",x"51",x"12",x"4a"),
   743 => (x"51",x"12",x"4a",x"a3"),
   744 => (x"12",x"4a",x"a3",x"d0"),
   745 => (x"4a",x"a3",x"d2",x"51"),
   746 => (x"a3",x"d4",x"51",x"12"),
   747 => (x"d6",x"51",x"12",x"4a"),
   748 => (x"51",x"12",x"4a",x"a3"),
   749 => (x"12",x"4a",x"a3",x"d8"),
   750 => (x"4a",x"a3",x"dc",x"51"),
   751 => (x"a3",x"de",x"51",x"12"),
   752 => (x"c1",x"51",x"12",x"4a"),
   753 => (x"87",x"fa",x"c0",x"7e"),
   754 => (x"99",x"c8",x"49",x"74"),
   755 => (x"87",x"eb",x"c0",x"05"),
   756 => (x"99",x"d0",x"49",x"74"),
   757 => (x"dc",x"87",x"d1",x"05"),
   758 => (x"cb",x"c0",x"02",x"66"),
   759 => (x"dc",x"49",x"73",x"87"),
   760 => (x"98",x"70",x"0f",x"66"),
   761 => (x"87",x"d3",x"c0",x"02"),
   762 => (x"c6",x"c0",x"05",x"6e"),
   763 => (x"ca",x"e5",x"c2",x"87"),
   764 => (x"c0",x"50",x"c0",x"48"),
   765 => (x"48",x"bf",x"e1",x"f2"),
   766 => (x"c2",x"87",x"e1",x"c2"),
   767 => (x"c0",x"48",x"d7",x"e5"),
   768 => (x"e5",x"c2",x"7e",x"50"),
   769 => (x"c2",x"49",x"bf",x"c6"),
   770 => (x"4a",x"bf",x"f6",x"dc"),
   771 => (x"fb",x"04",x"aa",x"71"),
   772 => (x"e9",x"c2",x"87",x"f7"),
   773 => (x"c0",x"05",x"bf",x"e7"),
   774 => (x"e5",x"c2",x"87",x"c8"),
   775 => (x"c1",x"02",x"bf",x"c2"),
   776 => (x"dc",x"c2",x"87",x"f8"),
   777 => (x"ed",x"49",x"bf",x"f2"),
   778 => (x"49",x"70",x"87",x"e4"),
   779 => (x"59",x"f6",x"dc",x"c2"),
   780 => (x"c2",x"48",x"a6",x"c4"),
   781 => (x"78",x"bf",x"f2",x"dc"),
   782 => (x"bf",x"c2",x"e5",x"c2"),
   783 => (x"87",x"d8",x"c0",x"02"),
   784 => (x"cf",x"49",x"66",x"c4"),
   785 => (x"f8",x"ff",x"ff",x"ff"),
   786 => (x"c0",x"02",x"a9",x"99"),
   787 => (x"4c",x"c0",x"87",x"c5"),
   788 => (x"c1",x"87",x"e1",x"c0"),
   789 => (x"87",x"dc",x"c0",x"4c"),
   790 => (x"cf",x"49",x"66",x"c4"),
   791 => (x"a9",x"99",x"f8",x"ff"),
   792 => (x"87",x"c8",x"c0",x"02"),
   793 => (x"c0",x"48",x"a6",x"c8"),
   794 => (x"87",x"c5",x"c0",x"78"),
   795 => (x"c1",x"48",x"a6",x"c8"),
   796 => (x"4c",x"66",x"c8",x"78"),
   797 => (x"c0",x"05",x"9c",x"74"),
   798 => (x"66",x"c4",x"87",x"e0"),
   799 => (x"c2",x"89",x"c2",x"49"),
   800 => (x"4a",x"bf",x"fa",x"e4"),
   801 => (x"d3",x"e9",x"c2",x"91"),
   802 => (x"dc",x"c2",x"4a",x"bf"),
   803 => (x"a1",x"72",x"48",x"ee"),
   804 => (x"f6",x"dc",x"c2",x"78"),
   805 => (x"f9",x"78",x"c0",x"48"),
   806 => (x"48",x"c0",x"87",x"df"),
   807 => (x"e5",x"eb",x"8e",x"f4"),
   808 => (x"00",x"00",x"00",x"87"),
   809 => (x"ff",x"ff",x"ff",x"00"),
   810 => (x"00",x"0c",x"b1",x"ff"),
   811 => (x"00",x"0c",x"ba",x"00"),
   812 => (x"54",x"41",x"46",x"00"),
   813 => (x"20",x"20",x"32",x"33"),
   814 => (x"41",x"46",x"00",x"20"),
   815 => (x"20",x"36",x"31",x"54"),
   816 => (x"1e",x"00",x"20",x"20"),
   817 => (x"c3",x"48",x"d4",x"ff"),
   818 => (x"48",x"68",x"78",x"ff"),
   819 => (x"ff",x"1e",x"4f",x"26"),
   820 => (x"ff",x"c3",x"48",x"d4"),
   821 => (x"48",x"d0",x"ff",x"78"),
   822 => (x"ff",x"78",x"e1",x"c0"),
   823 => (x"78",x"d4",x"48",x"d4"),
   824 => (x"48",x"eb",x"e9",x"c2"),
   825 => (x"50",x"bf",x"d4",x"ff"),
   826 => (x"ff",x"1e",x"4f",x"26"),
   827 => (x"e0",x"c0",x"48",x"d0"),
   828 => (x"1e",x"4f",x"26",x"78"),
   829 => (x"70",x"87",x"cc",x"ff"),
   830 => (x"c6",x"02",x"99",x"49"),
   831 => (x"a9",x"fb",x"c0",x"87"),
   832 => (x"71",x"87",x"f1",x"05"),
   833 => (x"0e",x"4f",x"26",x"48"),
   834 => (x"0e",x"5c",x"5b",x"5e"),
   835 => (x"4c",x"c0",x"4b",x"71"),
   836 => (x"70",x"87",x"f0",x"fe"),
   837 => (x"c0",x"02",x"99",x"49"),
   838 => (x"ec",x"c0",x"87",x"f9"),
   839 => (x"f2",x"c0",x"02",x"a9"),
   840 => (x"a9",x"fb",x"c0",x"87"),
   841 => (x"87",x"eb",x"c0",x"02"),
   842 => (x"ac",x"b7",x"66",x"cc"),
   843 => (x"d0",x"87",x"c7",x"03"),
   844 => (x"87",x"c2",x"02",x"66"),
   845 => (x"99",x"71",x"53",x"71"),
   846 => (x"c1",x"87",x"c2",x"02"),
   847 => (x"87",x"c3",x"fe",x"84"),
   848 => (x"02",x"99",x"49",x"70"),
   849 => (x"ec",x"c0",x"87",x"cd"),
   850 => (x"87",x"c7",x"02",x"a9"),
   851 => (x"05",x"a9",x"fb",x"c0"),
   852 => (x"d0",x"87",x"d5",x"ff"),
   853 => (x"87",x"c3",x"02",x"66"),
   854 => (x"c0",x"7b",x"97",x"c0"),
   855 => (x"c4",x"05",x"a9",x"ec"),
   856 => (x"c5",x"4a",x"74",x"87"),
   857 => (x"c0",x"4a",x"74",x"87"),
   858 => (x"48",x"72",x"8a",x"0a"),
   859 => (x"4d",x"26",x"87",x"c2"),
   860 => (x"4b",x"26",x"4c",x"26"),
   861 => (x"fd",x"1e",x"4f",x"26"),
   862 => (x"49",x"70",x"87",x"c9"),
   863 => (x"aa",x"f0",x"c0",x"4a"),
   864 => (x"c0",x"87",x"c9",x"04"),
   865 => (x"c3",x"01",x"aa",x"f9"),
   866 => (x"8a",x"f0",x"c0",x"87"),
   867 => (x"04",x"aa",x"c1",x"c1"),
   868 => (x"da",x"c1",x"87",x"c9"),
   869 => (x"87",x"c3",x"01",x"aa"),
   870 => (x"72",x"8a",x"f7",x"c0"),
   871 => (x"0e",x"4f",x"26",x"48"),
   872 => (x"0e",x"5c",x"5b",x"5e"),
   873 => (x"d4",x"ff",x"4a",x"71"),
   874 => (x"c0",x"49",x"72",x"4b"),
   875 => (x"4c",x"70",x"87",x"e7"),
   876 => (x"87",x"c2",x"02",x"9c"),
   877 => (x"d0",x"ff",x"8c",x"c1"),
   878 => (x"c1",x"78",x"c5",x"48"),
   879 => (x"49",x"74",x"7b",x"d5"),
   880 => (x"e5",x"c1",x"31",x"c6"),
   881 => (x"4a",x"bf",x"97",x"c8"),
   882 => (x"70",x"b0",x"71",x"48"),
   883 => (x"48",x"d0",x"ff",x"7b"),
   884 => (x"db",x"fe",x"78",x"c4"),
   885 => (x"5b",x"5e",x"0e",x"87"),
   886 => (x"f8",x"0e",x"5d",x"5c"),
   887 => (x"c0",x"4c",x"71",x"86"),
   888 => (x"87",x"ea",x"fb",x"7e"),
   889 => (x"fa",x"c0",x"4b",x"c0"),
   890 => (x"49",x"bf",x"97",x"c2"),
   891 => (x"cf",x"04",x"a9",x"c0"),
   892 => (x"87",x"ff",x"fb",x"87"),
   893 => (x"fa",x"c0",x"83",x"c1"),
   894 => (x"49",x"bf",x"97",x"c2"),
   895 => (x"87",x"f1",x"06",x"ab"),
   896 => (x"97",x"c2",x"fa",x"c0"),
   897 => (x"87",x"cf",x"02",x"bf"),
   898 => (x"70",x"87",x"f8",x"fa"),
   899 => (x"c6",x"02",x"99",x"49"),
   900 => (x"a9",x"ec",x"c0",x"87"),
   901 => (x"c0",x"87",x"f1",x"05"),
   902 => (x"87",x"e7",x"fa",x"4b"),
   903 => (x"e2",x"fa",x"4d",x"70"),
   904 => (x"58",x"a6",x"c8",x"87"),
   905 => (x"70",x"87",x"dc",x"fa"),
   906 => (x"c8",x"83",x"c1",x"4a"),
   907 => (x"69",x"97",x"49",x"a4"),
   908 => (x"c7",x"02",x"ad",x"49"),
   909 => (x"ad",x"ff",x"c0",x"87"),
   910 => (x"87",x"e7",x"c0",x"05"),
   911 => (x"97",x"49",x"a4",x"c9"),
   912 => (x"66",x"c4",x"49",x"69"),
   913 => (x"87",x"c7",x"02",x"a9"),
   914 => (x"a8",x"ff",x"c0",x"48"),
   915 => (x"ca",x"87",x"d4",x"05"),
   916 => (x"69",x"97",x"49",x"a4"),
   917 => (x"c6",x"02",x"aa",x"49"),
   918 => (x"aa",x"ff",x"c0",x"87"),
   919 => (x"c1",x"87",x"c4",x"05"),
   920 => (x"c0",x"87",x"d0",x"7e"),
   921 => (x"c6",x"02",x"ad",x"ec"),
   922 => (x"ad",x"fb",x"c0",x"87"),
   923 => (x"c0",x"87",x"c4",x"05"),
   924 => (x"6e",x"7e",x"c1",x"4b"),
   925 => (x"87",x"e1",x"fe",x"02"),
   926 => (x"73",x"87",x"ef",x"f9"),
   927 => (x"fb",x"8e",x"f8",x"48"),
   928 => (x"0e",x"00",x"87",x"ec"),
   929 => (x"5d",x"5c",x"5b",x"5e"),
   930 => (x"71",x"86",x"f8",x"0e"),
   931 => (x"4b",x"d4",x"ff",x"4d"),
   932 => (x"e9",x"c2",x"1e",x"75"),
   933 => (x"e7",x"e5",x"49",x"f0"),
   934 => (x"70",x"86",x"c4",x"87"),
   935 => (x"cc",x"c4",x"02",x"98"),
   936 => (x"48",x"a6",x"c4",x"87"),
   937 => (x"bf",x"ca",x"e5",x"c1"),
   938 => (x"fb",x"49",x"75",x"78"),
   939 => (x"d0",x"ff",x"87",x"f1"),
   940 => (x"c1",x"78",x"c5",x"48"),
   941 => (x"4a",x"c0",x"7b",x"d6"),
   942 => (x"11",x"49",x"a2",x"75"),
   943 => (x"cb",x"82",x"c1",x"7b"),
   944 => (x"f3",x"04",x"aa",x"b7"),
   945 => (x"c3",x"4a",x"cc",x"87"),
   946 => (x"82",x"c1",x"7b",x"ff"),
   947 => (x"aa",x"b7",x"e0",x"c0"),
   948 => (x"ff",x"87",x"f4",x"04"),
   949 => (x"78",x"c4",x"48",x"d0"),
   950 => (x"c5",x"7b",x"ff",x"c3"),
   951 => (x"7b",x"d3",x"c1",x"78"),
   952 => (x"78",x"c4",x"7b",x"c1"),
   953 => (x"b7",x"c0",x"48",x"66"),
   954 => (x"f0",x"c2",x"06",x"a8"),
   955 => (x"f8",x"e9",x"c2",x"87"),
   956 => (x"66",x"c4",x"4c",x"bf"),
   957 => (x"c8",x"88",x"74",x"48"),
   958 => (x"9c",x"74",x"58",x"a6"),
   959 => (x"87",x"f9",x"c1",x"02"),
   960 => (x"7e",x"fa",x"dc",x"c2"),
   961 => (x"8c",x"4d",x"c0",x"c8"),
   962 => (x"03",x"ac",x"b7",x"c0"),
   963 => (x"c0",x"c8",x"87",x"c6"),
   964 => (x"4c",x"c0",x"4d",x"a4"),
   965 => (x"97",x"eb",x"e9",x"c2"),
   966 => (x"99",x"d0",x"49",x"bf"),
   967 => (x"c0",x"87",x"d1",x"02"),
   968 => (x"f0",x"e9",x"c2",x"1e"),
   969 => (x"87",x"cc",x"e8",x"49"),
   970 => (x"49",x"70",x"86",x"c4"),
   971 => (x"87",x"ee",x"c0",x"4a"),
   972 => (x"1e",x"fa",x"dc",x"c2"),
   973 => (x"49",x"f0",x"e9",x"c2"),
   974 => (x"c4",x"87",x"f9",x"e7"),
   975 => (x"4a",x"49",x"70",x"86"),
   976 => (x"c8",x"48",x"d0",x"ff"),
   977 => (x"d4",x"c1",x"78",x"c5"),
   978 => (x"bf",x"97",x"6e",x"7b"),
   979 => (x"c1",x"48",x"6e",x"7b"),
   980 => (x"c1",x"7e",x"70",x"80"),
   981 => (x"f0",x"ff",x"05",x"8d"),
   982 => (x"48",x"d0",x"ff",x"87"),
   983 => (x"9a",x"72",x"78",x"c4"),
   984 => (x"c0",x"87",x"c5",x"05"),
   985 => (x"87",x"c7",x"c1",x"48"),
   986 => (x"e9",x"c2",x"1e",x"c1"),
   987 => (x"e9",x"e5",x"49",x"f0"),
   988 => (x"74",x"86",x"c4",x"87"),
   989 => (x"c7",x"fe",x"05",x"9c"),
   990 => (x"48",x"66",x"c4",x"87"),
   991 => (x"06",x"a8",x"b7",x"c0"),
   992 => (x"e9",x"c2",x"87",x"d1"),
   993 => (x"78",x"c0",x"48",x"f0"),
   994 => (x"78",x"c0",x"80",x"d0"),
   995 => (x"e9",x"c2",x"80",x"f4"),
   996 => (x"c4",x"78",x"bf",x"fc"),
   997 => (x"b7",x"c0",x"48",x"66"),
   998 => (x"d0",x"fd",x"01",x"a8"),
   999 => (x"48",x"d0",x"ff",x"87"),
  1000 => (x"d3",x"c1",x"78",x"c5"),
  1001 => (x"c4",x"7b",x"c0",x"7b"),
  1002 => (x"c2",x"48",x"c1",x"78"),
  1003 => (x"f8",x"48",x"c0",x"87"),
  1004 => (x"26",x"4d",x"26",x"8e"),
  1005 => (x"26",x"4b",x"26",x"4c"),
  1006 => (x"5b",x"5e",x"0e",x"4f"),
  1007 => (x"1e",x"0e",x"5d",x"5c"),
  1008 => (x"4c",x"c0",x"4b",x"71"),
  1009 => (x"c0",x"04",x"ab",x"4d"),
  1010 => (x"f7",x"c0",x"87",x"e8"),
  1011 => (x"9d",x"75",x"1e",x"d5"),
  1012 => (x"c0",x"87",x"c4",x"02"),
  1013 => (x"c1",x"87",x"c2",x"4a"),
  1014 => (x"eb",x"49",x"72",x"4a"),
  1015 => (x"86",x"c4",x"87",x"ec"),
  1016 => (x"84",x"c1",x"7e",x"70"),
  1017 => (x"87",x"c2",x"05",x"6e"),
  1018 => (x"85",x"c1",x"4c",x"73"),
  1019 => (x"ff",x"06",x"ac",x"73"),
  1020 => (x"48",x"6e",x"87",x"d8"),
  1021 => (x"87",x"f9",x"fe",x"26"),
  1022 => (x"5c",x"5b",x"5e",x"0e"),
  1023 => (x"cc",x"4b",x"71",x"0e"),
  1024 => (x"87",x"d8",x"02",x"66"),
  1025 => (x"8c",x"f0",x"c0",x"4c"),
  1026 => (x"74",x"87",x"d8",x"02"),
  1027 => (x"02",x"8a",x"c1",x"4a"),
  1028 => (x"02",x"8a",x"87",x"d1"),
  1029 => (x"02",x"8a",x"87",x"cd"),
  1030 => (x"87",x"d9",x"87",x"c9"),
  1031 => (x"e2",x"f9",x"49",x"73"),
  1032 => (x"74",x"87",x"d2",x"87"),
  1033 => (x"c1",x"49",x"c0",x"1e"),
  1034 => (x"74",x"87",x"e6",x"d9"),
  1035 => (x"c1",x"49",x"73",x"1e"),
  1036 => (x"c8",x"87",x"de",x"d9"),
  1037 => (x"87",x"fb",x"fd",x"86"),
  1038 => (x"5c",x"5b",x"5e",x"0e"),
  1039 => (x"71",x"1e",x"0e",x"5d"),
  1040 => (x"91",x"de",x"49",x"4c"),
  1041 => (x"4d",x"d8",x"ea",x"c2"),
  1042 => (x"6d",x"97",x"85",x"71"),
  1043 => (x"87",x"dd",x"c1",x"02"),
  1044 => (x"bf",x"c4",x"ea",x"c2"),
  1045 => (x"72",x"82",x"74",x"4a"),
  1046 => (x"87",x"dd",x"fd",x"49"),
  1047 => (x"98",x"48",x"7e",x"70"),
  1048 => (x"87",x"f2",x"c0",x"02"),
  1049 => (x"4b",x"cc",x"ea",x"c2"),
  1050 => (x"49",x"cb",x"4a",x"70"),
  1051 => (x"87",x"f7",x"c0",x"ff"),
  1052 => (x"93",x"cb",x"4b",x"74"),
  1053 => (x"83",x"dc",x"e5",x"c1"),
  1054 => (x"c2",x"c1",x"83",x"c4"),
  1055 => (x"49",x"74",x"7b",x"f1"),
  1056 => (x"87",x"f9",x"c2",x"c1"),
  1057 => (x"e5",x"c1",x"7b",x"75"),
  1058 => (x"49",x"bf",x"97",x"c9"),
  1059 => (x"cc",x"ea",x"c2",x"1e"),
  1060 => (x"87",x"e4",x"fd",x"49"),
  1061 => (x"49",x"74",x"86",x"c4"),
  1062 => (x"87",x"e1",x"c2",x"c1"),
  1063 => (x"c4",x"c1",x"49",x"c0"),
  1064 => (x"e9",x"c2",x"87",x"c0"),
  1065 => (x"78",x"c0",x"48",x"ec"),
  1066 => (x"de",x"de",x"49",x"c1"),
  1067 => (x"c0",x"fc",x"26",x"87"),
  1068 => (x"61",x"6f",x"4c",x"87"),
  1069 => (x"67",x"6e",x"69",x"64"),
  1070 => (x"00",x"2e",x"2e",x"2e"),
  1071 => (x"5c",x"5b",x"5e",x"0e"),
  1072 => (x"4a",x"4b",x"71",x"0e"),
  1073 => (x"bf",x"c4",x"ea",x"c2"),
  1074 => (x"fb",x"49",x"72",x"82"),
  1075 => (x"4c",x"70",x"87",x"eb"),
  1076 => (x"87",x"c4",x"02",x"9c"),
  1077 => (x"87",x"fa",x"e6",x"49"),
  1078 => (x"48",x"c4",x"ea",x"c2"),
  1079 => (x"49",x"c1",x"78",x"c0"),
  1080 => (x"fb",x"87",x"e8",x"dd"),
  1081 => (x"5e",x"0e",x"87",x"cd"),
  1082 => (x"0e",x"5d",x"5c",x"5b"),
  1083 => (x"dc",x"c2",x"86",x"f4"),
  1084 => (x"4c",x"c0",x"4d",x"fa"),
  1085 => (x"c0",x"48",x"a6",x"c4"),
  1086 => (x"c4",x"ea",x"c2",x"78"),
  1087 => (x"a9",x"c0",x"49",x"bf"),
  1088 => (x"87",x"c1",x"c1",x"06"),
  1089 => (x"48",x"fa",x"dc",x"c2"),
  1090 => (x"f8",x"c0",x"02",x"98"),
  1091 => (x"d5",x"f7",x"c0",x"87"),
  1092 => (x"02",x"66",x"c8",x"1e"),
  1093 => (x"a6",x"c4",x"87",x"c7"),
  1094 => (x"c5",x"78",x"c0",x"48"),
  1095 => (x"48",x"a6",x"c4",x"87"),
  1096 => (x"66",x"c4",x"78",x"c1"),
  1097 => (x"87",x"e2",x"e6",x"49"),
  1098 => (x"4d",x"70",x"86",x"c4"),
  1099 => (x"66",x"c4",x"84",x"c1"),
  1100 => (x"c8",x"80",x"c1",x"48"),
  1101 => (x"ea",x"c2",x"58",x"a6"),
  1102 => (x"ac",x"49",x"bf",x"c4"),
  1103 => (x"75",x"87",x"c6",x"03"),
  1104 => (x"c8",x"ff",x"05",x"9d"),
  1105 => (x"75",x"4c",x"c0",x"87"),
  1106 => (x"e0",x"c3",x"02",x"9d"),
  1107 => (x"d5",x"f7",x"c0",x"87"),
  1108 => (x"02",x"66",x"c8",x"1e"),
  1109 => (x"a6",x"cc",x"87",x"c7"),
  1110 => (x"c5",x"78",x"c0",x"48"),
  1111 => (x"48",x"a6",x"cc",x"87"),
  1112 => (x"66",x"cc",x"78",x"c1"),
  1113 => (x"87",x"e2",x"e5",x"49"),
  1114 => (x"7e",x"70",x"86",x"c4"),
  1115 => (x"c2",x"02",x"98",x"48"),
  1116 => (x"cb",x"49",x"87",x"e8"),
  1117 => (x"49",x"69",x"97",x"81"),
  1118 => (x"c1",x"02",x"99",x"d0"),
  1119 => (x"c2",x"c1",x"87",x"d6"),
  1120 => (x"49",x"74",x"4a",x"fc"),
  1121 => (x"e5",x"c1",x"91",x"cb"),
  1122 => (x"79",x"72",x"81",x"dc"),
  1123 => (x"ff",x"c3",x"81",x"c8"),
  1124 => (x"de",x"49",x"74",x"51"),
  1125 => (x"d8",x"ea",x"c2",x"91"),
  1126 => (x"c2",x"85",x"71",x"4d"),
  1127 => (x"c1",x"7d",x"97",x"c1"),
  1128 => (x"e0",x"c0",x"49",x"a5"),
  1129 => (x"ca",x"e5",x"c2",x"51"),
  1130 => (x"d2",x"02",x"bf",x"97"),
  1131 => (x"c2",x"84",x"c1",x"87"),
  1132 => (x"e5",x"c2",x"4b",x"a5"),
  1133 => (x"49",x"db",x"4a",x"ca"),
  1134 => (x"87",x"eb",x"fb",x"fe"),
  1135 => (x"cd",x"87",x"db",x"c1"),
  1136 => (x"51",x"c0",x"49",x"a5"),
  1137 => (x"a5",x"c2",x"84",x"c1"),
  1138 => (x"cb",x"4a",x"6e",x"4b"),
  1139 => (x"d6",x"fb",x"fe",x"49"),
  1140 => (x"87",x"c6",x"c1",x"87"),
  1141 => (x"4a",x"f8",x"c0",x"c1"),
  1142 => (x"91",x"cb",x"49",x"74"),
  1143 => (x"81",x"dc",x"e5",x"c1"),
  1144 => (x"e5",x"c2",x"79",x"72"),
  1145 => (x"02",x"bf",x"97",x"ca"),
  1146 => (x"49",x"74",x"87",x"d8"),
  1147 => (x"84",x"c1",x"91",x"de"),
  1148 => (x"4b",x"d8",x"ea",x"c2"),
  1149 => (x"e5",x"c2",x"83",x"71"),
  1150 => (x"49",x"dd",x"4a",x"ca"),
  1151 => (x"87",x"e7",x"fa",x"fe"),
  1152 => (x"4b",x"74",x"87",x"d8"),
  1153 => (x"ea",x"c2",x"93",x"de"),
  1154 => (x"a3",x"cb",x"83",x"d8"),
  1155 => (x"c1",x"51",x"c0",x"49"),
  1156 => (x"4a",x"6e",x"73",x"84"),
  1157 => (x"fa",x"fe",x"49",x"cb"),
  1158 => (x"66",x"c4",x"87",x"cd"),
  1159 => (x"c8",x"80",x"c1",x"48"),
  1160 => (x"ac",x"c7",x"58",x"a6"),
  1161 => (x"87",x"c5",x"c0",x"03"),
  1162 => (x"e0",x"fc",x"05",x"6e"),
  1163 => (x"f4",x"48",x"74",x"87"),
  1164 => (x"87",x"fd",x"f5",x"8e"),
  1165 => (x"71",x"1e",x"73",x"1e"),
  1166 => (x"91",x"cb",x"49",x"4b"),
  1167 => (x"81",x"dc",x"e5",x"c1"),
  1168 => (x"c1",x"4a",x"a1",x"c8"),
  1169 => (x"12",x"48",x"c8",x"e5"),
  1170 => (x"4a",x"a1",x"c9",x"50"),
  1171 => (x"48",x"c2",x"fa",x"c0"),
  1172 => (x"81",x"ca",x"50",x"12"),
  1173 => (x"48",x"c9",x"e5",x"c1"),
  1174 => (x"e5",x"c1",x"50",x"11"),
  1175 => (x"49",x"bf",x"97",x"c9"),
  1176 => (x"f6",x"49",x"c0",x"1e"),
  1177 => (x"e9",x"c2",x"87",x"d2"),
  1178 => (x"78",x"de",x"48",x"ec"),
  1179 => (x"da",x"d7",x"49",x"c1"),
  1180 => (x"c0",x"f5",x"26",x"87"),
  1181 => (x"4a",x"71",x"1e",x"87"),
  1182 => (x"c1",x"91",x"cb",x"49"),
  1183 => (x"c8",x"81",x"dc",x"e5"),
  1184 => (x"c2",x"48",x"11",x"81"),
  1185 => (x"c2",x"58",x"f0",x"e9"),
  1186 => (x"c0",x"48",x"c4",x"ea"),
  1187 => (x"d6",x"49",x"c1",x"78"),
  1188 => (x"4f",x"26",x"87",x"f9"),
  1189 => (x"c0",x"49",x"c0",x"1e"),
  1190 => (x"26",x"87",x"c7",x"fc"),
  1191 => (x"99",x"71",x"1e",x"4f"),
  1192 => (x"c1",x"87",x"d2",x"02"),
  1193 => (x"c0",x"48",x"f1",x"e6"),
  1194 => (x"c1",x"80",x"f7",x"50"),
  1195 => (x"c1",x"40",x"f5",x"c9"),
  1196 => (x"ce",x"78",x"d5",x"e5"),
  1197 => (x"ed",x"e6",x"c1",x"87"),
  1198 => (x"ce",x"e5",x"c1",x"48"),
  1199 => (x"c1",x"80",x"fc",x"78"),
  1200 => (x"26",x"78",x"d4",x"ca"),
  1201 => (x"5b",x"5e",x"0e",x"4f"),
  1202 => (x"f4",x"0e",x"5d",x"5c"),
  1203 => (x"49",x"4d",x"71",x"86"),
  1204 => (x"e5",x"c1",x"91",x"cb"),
  1205 => (x"a1",x"c8",x"81",x"dc"),
  1206 => (x"7e",x"a1",x"ca",x"4a"),
  1207 => (x"c2",x"48",x"a6",x"c4"),
  1208 => (x"78",x"bf",x"f4",x"ed"),
  1209 => (x"4b",x"bf",x"97",x"6e"),
  1210 => (x"73",x"48",x"66",x"c4"),
  1211 => (x"4c",x"4b",x"70",x"28"),
  1212 => (x"a6",x"cc",x"48",x"12"),
  1213 => (x"c1",x"9c",x"70",x"58"),
  1214 => (x"97",x"81",x"c9",x"84"),
  1215 => (x"ac",x"b7",x"49",x"69"),
  1216 => (x"c0",x"87",x"c2",x"04"),
  1217 => (x"bf",x"97",x"6e",x"4c"),
  1218 => (x"49",x"66",x"c8",x"4a"),
  1219 => (x"b9",x"ff",x"31",x"72"),
  1220 => (x"74",x"99",x"66",x"c4"),
  1221 => (x"70",x"30",x"72",x"48"),
  1222 => (x"b0",x"71",x"48",x"4a"),
  1223 => (x"58",x"f8",x"ed",x"c2"),
  1224 => (x"87",x"d9",x"e6",x"c0"),
  1225 => (x"e2",x"d4",x"49",x"c0"),
  1226 => (x"c0",x"49",x"75",x"87"),
  1227 => (x"f4",x"87",x"ce",x"f8"),
  1228 => (x"87",x"fd",x"f1",x"8e"),
  1229 => (x"71",x"1e",x"73",x"1e"),
  1230 => (x"c8",x"fe",x"49",x"4b"),
  1231 => (x"fe",x"49",x"73",x"87"),
  1232 => (x"f0",x"f1",x"87",x"c3"),
  1233 => (x"1e",x"73",x"1e",x"87"),
  1234 => (x"a3",x"c6",x"4b",x"71"),
  1235 => (x"87",x"db",x"02",x"4a"),
  1236 => (x"d6",x"02",x"8a",x"c1"),
  1237 => (x"c1",x"02",x"8a",x"87"),
  1238 => (x"02",x"8a",x"87",x"da"),
  1239 => (x"8a",x"87",x"fc",x"c0"),
  1240 => (x"87",x"e1",x"c0",x"02"),
  1241 => (x"87",x"cb",x"02",x"8a"),
  1242 => (x"c7",x"87",x"db",x"c1"),
  1243 => (x"87",x"c5",x"fc",x"49"),
  1244 => (x"c2",x"87",x"de",x"c1"),
  1245 => (x"02",x"bf",x"c4",x"ea"),
  1246 => (x"48",x"87",x"cb",x"c1"),
  1247 => (x"ea",x"c2",x"88",x"c1"),
  1248 => (x"c1",x"c1",x"58",x"c8"),
  1249 => (x"c8",x"ea",x"c2",x"87"),
  1250 => (x"f9",x"c0",x"02",x"bf"),
  1251 => (x"c4",x"ea",x"c2",x"87"),
  1252 => (x"80",x"c1",x"48",x"bf"),
  1253 => (x"58",x"c8",x"ea",x"c2"),
  1254 => (x"c2",x"87",x"eb",x"c0"),
  1255 => (x"49",x"bf",x"c4",x"ea"),
  1256 => (x"ea",x"c2",x"89",x"c6"),
  1257 => (x"b7",x"c0",x"59",x"c8"),
  1258 => (x"87",x"da",x"03",x"a9"),
  1259 => (x"48",x"c4",x"ea",x"c2"),
  1260 => (x"87",x"d2",x"78",x"c0"),
  1261 => (x"bf",x"c8",x"ea",x"c2"),
  1262 => (x"c2",x"87",x"cb",x"02"),
  1263 => (x"48",x"bf",x"c4",x"ea"),
  1264 => (x"ea",x"c2",x"80",x"c6"),
  1265 => (x"49",x"c0",x"58",x"c8"),
  1266 => (x"73",x"87",x"c0",x"d2"),
  1267 => (x"ec",x"f5",x"c0",x"49"),
  1268 => (x"87",x"e1",x"ef",x"87"),
  1269 => (x"5c",x"5b",x"5e",x"0e"),
  1270 => (x"d0",x"ff",x"0e",x"5d"),
  1271 => (x"59",x"a6",x"dc",x"86"),
  1272 => (x"c0",x"48",x"a6",x"c8"),
  1273 => (x"c1",x"80",x"c4",x"78"),
  1274 => (x"c4",x"78",x"66",x"c4"),
  1275 => (x"c4",x"78",x"c1",x"80"),
  1276 => (x"c2",x"78",x"c1",x"80"),
  1277 => (x"c1",x"48",x"c8",x"ea"),
  1278 => (x"ec",x"e9",x"c2",x"78"),
  1279 => (x"a8",x"de",x"48",x"bf"),
  1280 => (x"f3",x"87",x"cb",x"05"),
  1281 => (x"49",x"70",x"87",x"e0"),
  1282 => (x"cf",x"59",x"a6",x"cc"),
  1283 => (x"fd",x"e2",x"87",x"fc"),
  1284 => (x"87",x"df",x"e3",x"87"),
  1285 => (x"70",x"87",x"ec",x"e2"),
  1286 => (x"ac",x"fb",x"c0",x"4c"),
  1287 => (x"87",x"fb",x"c1",x"02"),
  1288 => (x"c1",x"05",x"66",x"d8"),
  1289 => (x"c0",x"c1",x"87",x"ed"),
  1290 => (x"82",x"c4",x"4a",x"66"),
  1291 => (x"1e",x"72",x"7e",x"6a"),
  1292 => (x"48",x"ff",x"e0",x"c1"),
  1293 => (x"c8",x"49",x"66",x"c4"),
  1294 => (x"41",x"20",x"4a",x"a1"),
  1295 => (x"f9",x"05",x"aa",x"71"),
  1296 => (x"26",x"51",x"10",x"87"),
  1297 => (x"66",x"c0",x"c1",x"4a"),
  1298 => (x"f4",x"c8",x"c1",x"48"),
  1299 => (x"c7",x"49",x"6a",x"78"),
  1300 => (x"c1",x"51",x"74",x"81"),
  1301 => (x"c8",x"49",x"66",x"c0"),
  1302 => (x"c1",x"51",x"c1",x"81"),
  1303 => (x"c9",x"49",x"66",x"c0"),
  1304 => (x"c1",x"51",x"c0",x"81"),
  1305 => (x"ca",x"49",x"66",x"c0"),
  1306 => (x"c1",x"51",x"c0",x"81"),
  1307 => (x"6a",x"1e",x"d8",x"1e"),
  1308 => (x"e2",x"81",x"c8",x"49"),
  1309 => (x"86",x"c8",x"87",x"d1"),
  1310 => (x"48",x"66",x"c4",x"c1"),
  1311 => (x"c7",x"01",x"a8",x"c0"),
  1312 => (x"48",x"a6",x"c8",x"87"),
  1313 => (x"87",x"ce",x"78",x"c1"),
  1314 => (x"48",x"66",x"c4",x"c1"),
  1315 => (x"a6",x"d0",x"88",x"c1"),
  1316 => (x"e1",x"87",x"c3",x"58"),
  1317 => (x"a6",x"d0",x"87",x"dd"),
  1318 => (x"74",x"78",x"c2",x"48"),
  1319 => (x"e5",x"cd",x"02",x"9c"),
  1320 => (x"48",x"66",x"c8",x"87"),
  1321 => (x"a8",x"66",x"c8",x"c1"),
  1322 => (x"87",x"da",x"cd",x"03"),
  1323 => (x"c0",x"48",x"a6",x"dc"),
  1324 => (x"c0",x"80",x"e8",x"78"),
  1325 => (x"87",x"cb",x"e0",x"78"),
  1326 => (x"d0",x"c1",x"4c",x"70"),
  1327 => (x"da",x"c2",x"05",x"ac"),
  1328 => (x"7e",x"66",x"c4",x"87"),
  1329 => (x"70",x"87",x"ef",x"e2"),
  1330 => (x"59",x"a6",x"c8",x"49"),
  1331 => (x"87",x"f3",x"df",x"ff"),
  1332 => (x"ec",x"c0",x"4c",x"70"),
  1333 => (x"ed",x"c1",x"05",x"ac"),
  1334 => (x"49",x"66",x"c8",x"87"),
  1335 => (x"c0",x"c1",x"91",x"cb"),
  1336 => (x"a1",x"c4",x"81",x"66"),
  1337 => (x"c8",x"4d",x"6a",x"4a"),
  1338 => (x"66",x"c4",x"4a",x"a1"),
  1339 => (x"f5",x"c9",x"c1",x"52"),
  1340 => (x"ce",x"df",x"ff",x"79"),
  1341 => (x"9c",x"4c",x"70",x"87"),
  1342 => (x"c0",x"87",x"d9",x"02"),
  1343 => (x"d3",x"02",x"ac",x"fb"),
  1344 => (x"ff",x"55",x"74",x"87"),
  1345 => (x"70",x"87",x"fc",x"de"),
  1346 => (x"c7",x"02",x"9c",x"4c"),
  1347 => (x"ac",x"fb",x"c0",x"87"),
  1348 => (x"87",x"ed",x"ff",x"05"),
  1349 => (x"c2",x"55",x"e0",x"c0"),
  1350 => (x"97",x"c0",x"55",x"c1"),
  1351 => (x"49",x"66",x"d8",x"7d"),
  1352 => (x"db",x"05",x"a9",x"6e"),
  1353 => (x"48",x"66",x"c8",x"87"),
  1354 => (x"04",x"a8",x"66",x"cc"),
  1355 => (x"66",x"c8",x"87",x"ca"),
  1356 => (x"cc",x"80",x"c1",x"48"),
  1357 => (x"87",x"c8",x"58",x"a6"),
  1358 => (x"c1",x"48",x"66",x"cc"),
  1359 => (x"58",x"a6",x"d0",x"88"),
  1360 => (x"87",x"ff",x"dd",x"ff"),
  1361 => (x"d0",x"c1",x"4c",x"70"),
  1362 => (x"87",x"c8",x"05",x"ac"),
  1363 => (x"c1",x"48",x"66",x"d4"),
  1364 => (x"58",x"a6",x"d8",x"80"),
  1365 => (x"02",x"ac",x"d0",x"c1"),
  1366 => (x"c0",x"87",x"e6",x"fd"),
  1367 => (x"d8",x"48",x"a6",x"e0"),
  1368 => (x"66",x"c4",x"78",x"66"),
  1369 => (x"66",x"e0",x"c0",x"48"),
  1370 => (x"eb",x"c9",x"05",x"a8"),
  1371 => (x"a6",x"e4",x"c0",x"87"),
  1372 => (x"74",x"78",x"c0",x"48"),
  1373 => (x"88",x"fb",x"c0",x"48"),
  1374 => (x"98",x"48",x"7e",x"70"),
  1375 => (x"87",x"ed",x"c9",x"02"),
  1376 => (x"70",x"88",x"cb",x"48"),
  1377 => (x"02",x"98",x"48",x"7e"),
  1378 => (x"48",x"87",x"cd",x"c1"),
  1379 => (x"7e",x"70",x"88",x"c9"),
  1380 => (x"c4",x"02",x"98",x"48"),
  1381 => (x"c4",x"48",x"87",x"c1"),
  1382 => (x"48",x"7e",x"70",x"88"),
  1383 => (x"87",x"ce",x"02",x"98"),
  1384 => (x"70",x"88",x"c1",x"48"),
  1385 => (x"02",x"98",x"48",x"7e"),
  1386 => (x"c8",x"87",x"ec",x"c3"),
  1387 => (x"a6",x"dc",x"87",x"e1"),
  1388 => (x"78",x"f0",x"c0",x"48"),
  1389 => (x"87",x"cb",x"dc",x"ff"),
  1390 => (x"ec",x"c0",x"4c",x"70"),
  1391 => (x"c4",x"c0",x"02",x"ac"),
  1392 => (x"a6",x"e0",x"c0",x"87"),
  1393 => (x"ac",x"ec",x"c0",x"5c"),
  1394 => (x"ff",x"87",x"cd",x"02"),
  1395 => (x"70",x"87",x"f4",x"db"),
  1396 => (x"ac",x"ec",x"c0",x"4c"),
  1397 => (x"87",x"f3",x"ff",x"05"),
  1398 => (x"02",x"ac",x"ec",x"c0"),
  1399 => (x"ff",x"87",x"c4",x"c0"),
  1400 => (x"c0",x"87",x"e0",x"db"),
  1401 => (x"d0",x"1e",x"ca",x"1e"),
  1402 => (x"91",x"cb",x"49",x"66"),
  1403 => (x"48",x"66",x"c8",x"c1"),
  1404 => (x"a6",x"cc",x"80",x"71"),
  1405 => (x"48",x"66",x"c8",x"58"),
  1406 => (x"a6",x"d0",x"80",x"c4"),
  1407 => (x"bf",x"66",x"cc",x"58"),
  1408 => (x"c2",x"dc",x"ff",x"49"),
  1409 => (x"de",x"1e",x"c1",x"87"),
  1410 => (x"bf",x"66",x"d4",x"1e"),
  1411 => (x"f6",x"db",x"ff",x"49"),
  1412 => (x"70",x"86",x"d0",x"87"),
  1413 => (x"89",x"09",x"c0",x"49"),
  1414 => (x"59",x"a6",x"ec",x"c0"),
  1415 => (x"48",x"66",x"e8",x"c0"),
  1416 => (x"c0",x"06",x"a8",x"c0"),
  1417 => (x"e8",x"c0",x"87",x"ee"),
  1418 => (x"a8",x"dd",x"48",x"66"),
  1419 => (x"87",x"e4",x"c0",x"03"),
  1420 => (x"49",x"bf",x"66",x"c4"),
  1421 => (x"81",x"66",x"e8",x"c0"),
  1422 => (x"c0",x"51",x"e0",x"c0"),
  1423 => (x"c1",x"49",x"66",x"e8"),
  1424 => (x"bf",x"66",x"c4",x"81"),
  1425 => (x"51",x"c1",x"c2",x"81"),
  1426 => (x"49",x"66",x"e8",x"c0"),
  1427 => (x"66",x"c4",x"81",x"c2"),
  1428 => (x"51",x"c0",x"81",x"bf"),
  1429 => (x"c8",x"c1",x"48",x"6e"),
  1430 => (x"49",x"6e",x"78",x"f4"),
  1431 => (x"66",x"d0",x"81",x"c8"),
  1432 => (x"c9",x"49",x"6e",x"51"),
  1433 => (x"51",x"66",x"d4",x"81"),
  1434 => (x"81",x"ca",x"49",x"6e"),
  1435 => (x"d0",x"51",x"66",x"dc"),
  1436 => (x"80",x"c1",x"48",x"66"),
  1437 => (x"c8",x"58",x"a6",x"d4"),
  1438 => (x"66",x"cc",x"48",x"66"),
  1439 => (x"cb",x"c0",x"04",x"a8"),
  1440 => (x"48",x"66",x"c8",x"87"),
  1441 => (x"a6",x"cc",x"80",x"c1"),
  1442 => (x"87",x"e1",x"c5",x"58"),
  1443 => (x"c1",x"48",x"66",x"cc"),
  1444 => (x"58",x"a6",x"d0",x"88"),
  1445 => (x"ff",x"87",x"d6",x"c5"),
  1446 => (x"70",x"87",x"db",x"db"),
  1447 => (x"a6",x"ec",x"c0",x"49"),
  1448 => (x"d1",x"db",x"ff",x"59"),
  1449 => (x"c0",x"49",x"70",x"87"),
  1450 => (x"dc",x"59",x"a6",x"e0"),
  1451 => (x"ec",x"c0",x"48",x"66"),
  1452 => (x"ca",x"c0",x"05",x"a8"),
  1453 => (x"48",x"a6",x"dc",x"87"),
  1454 => (x"78",x"66",x"e8",x"c0"),
  1455 => (x"ff",x"87",x"c4",x"c0"),
  1456 => (x"c8",x"87",x"c0",x"d8"),
  1457 => (x"91",x"cb",x"49",x"66"),
  1458 => (x"48",x"66",x"c0",x"c1"),
  1459 => (x"7e",x"70",x"80",x"71"),
  1460 => (x"6e",x"82",x"c8",x"4a"),
  1461 => (x"c0",x"81",x"ca",x"49"),
  1462 => (x"dc",x"51",x"66",x"e8"),
  1463 => (x"81",x"c1",x"49",x"66"),
  1464 => (x"89",x"66",x"e8",x"c0"),
  1465 => (x"30",x"71",x"48",x"c1"),
  1466 => (x"89",x"c1",x"49",x"70"),
  1467 => (x"c2",x"7a",x"97",x"71"),
  1468 => (x"49",x"bf",x"f4",x"ed"),
  1469 => (x"29",x"66",x"e8",x"c0"),
  1470 => (x"48",x"4a",x"6a",x"97"),
  1471 => (x"f0",x"c0",x"98",x"71"),
  1472 => (x"49",x"6e",x"58",x"a6"),
  1473 => (x"4d",x"69",x"81",x"c4"),
  1474 => (x"48",x"66",x"e0",x"c0"),
  1475 => (x"02",x"a8",x"66",x"c4"),
  1476 => (x"c4",x"87",x"c8",x"c0"),
  1477 => (x"78",x"c0",x"48",x"a6"),
  1478 => (x"c4",x"87",x"c5",x"c0"),
  1479 => (x"78",x"c1",x"48",x"a6"),
  1480 => (x"c0",x"1e",x"66",x"c4"),
  1481 => (x"49",x"75",x"1e",x"e0"),
  1482 => (x"87",x"db",x"d7",x"ff"),
  1483 => (x"4c",x"70",x"86",x"c8"),
  1484 => (x"06",x"ac",x"b7",x"c0"),
  1485 => (x"74",x"87",x"d4",x"c1"),
  1486 => (x"49",x"e0",x"c0",x"85"),
  1487 => (x"4b",x"75",x"89",x"74"),
  1488 => (x"4a",x"c8",x"e1",x"c1"),
  1489 => (x"de",x"e5",x"fe",x"71"),
  1490 => (x"c0",x"85",x"c2",x"87"),
  1491 => (x"c1",x"48",x"66",x"e4"),
  1492 => (x"a6",x"e8",x"c0",x"80"),
  1493 => (x"66",x"ec",x"c0",x"58"),
  1494 => (x"70",x"81",x"c1",x"49"),
  1495 => (x"c8",x"c0",x"02",x"a9"),
  1496 => (x"48",x"a6",x"c4",x"87"),
  1497 => (x"c5",x"c0",x"78",x"c0"),
  1498 => (x"48",x"a6",x"c4",x"87"),
  1499 => (x"66",x"c4",x"78",x"c1"),
  1500 => (x"49",x"a4",x"c2",x"1e"),
  1501 => (x"71",x"48",x"e0",x"c0"),
  1502 => (x"1e",x"49",x"70",x"88"),
  1503 => (x"d6",x"ff",x"49",x"75"),
  1504 => (x"86",x"c8",x"87",x"c5"),
  1505 => (x"01",x"a8",x"b7",x"c0"),
  1506 => (x"c0",x"87",x"c0",x"ff"),
  1507 => (x"c0",x"02",x"66",x"e4"),
  1508 => (x"49",x"6e",x"87",x"d1"),
  1509 => (x"e4",x"c0",x"81",x"c9"),
  1510 => (x"48",x"6e",x"51",x"66"),
  1511 => (x"78",x"c5",x"cb",x"c1"),
  1512 => (x"6e",x"87",x"cc",x"c0"),
  1513 => (x"c2",x"81",x"c9",x"49"),
  1514 => (x"c1",x"48",x"6e",x"51"),
  1515 => (x"c8",x"78",x"f4",x"cc"),
  1516 => (x"66",x"cc",x"48",x"66"),
  1517 => (x"cb",x"c0",x"04",x"a8"),
  1518 => (x"48",x"66",x"c8",x"87"),
  1519 => (x"a6",x"cc",x"80",x"c1"),
  1520 => (x"87",x"e9",x"c0",x"58"),
  1521 => (x"c1",x"48",x"66",x"cc"),
  1522 => (x"58",x"a6",x"d0",x"88"),
  1523 => (x"ff",x"87",x"de",x"c0"),
  1524 => (x"70",x"87",x"e0",x"d4"),
  1525 => (x"87",x"d5",x"c0",x"4c"),
  1526 => (x"05",x"ac",x"c6",x"c1"),
  1527 => (x"d0",x"87",x"c8",x"c0"),
  1528 => (x"80",x"c1",x"48",x"66"),
  1529 => (x"ff",x"58",x"a6",x"d4"),
  1530 => (x"70",x"87",x"c8",x"d4"),
  1531 => (x"48",x"66",x"d4",x"4c"),
  1532 => (x"a6",x"d8",x"80",x"c1"),
  1533 => (x"02",x"9c",x"74",x"58"),
  1534 => (x"c8",x"87",x"cb",x"c0"),
  1535 => (x"c8",x"c1",x"48",x"66"),
  1536 => (x"f2",x"04",x"a8",x"66"),
  1537 => (x"d3",x"ff",x"87",x"e6"),
  1538 => (x"66",x"c8",x"87",x"e0"),
  1539 => (x"03",x"a8",x"c7",x"48"),
  1540 => (x"c2",x"87",x"e5",x"c0"),
  1541 => (x"c0",x"48",x"c8",x"ea"),
  1542 => (x"49",x"66",x"c8",x"78"),
  1543 => (x"c0",x"c1",x"91",x"cb"),
  1544 => (x"a1",x"c4",x"81",x"66"),
  1545 => (x"c0",x"4a",x"6a",x"4a"),
  1546 => (x"66",x"c8",x"79",x"52"),
  1547 => (x"cc",x"80",x"c1",x"48"),
  1548 => (x"a8",x"c7",x"58",x"a6"),
  1549 => (x"87",x"db",x"ff",x"04"),
  1550 => (x"ff",x"8e",x"d0",x"ff"),
  1551 => (x"4c",x"87",x"f2",x"dd"),
  1552 => (x"20",x"64",x"61",x"6f"),
  1553 => (x"00",x"20",x"2e",x"2a"),
  1554 => (x"1e",x"00",x"20",x"3a"),
  1555 => (x"4b",x"71",x"1e",x"73"),
  1556 => (x"87",x"c6",x"02",x"9b"),
  1557 => (x"48",x"c4",x"ea",x"c2"),
  1558 => (x"1e",x"c7",x"78",x"c0"),
  1559 => (x"bf",x"c4",x"ea",x"c2"),
  1560 => (x"e5",x"c1",x"1e",x"49"),
  1561 => (x"e9",x"c2",x"1e",x"dc"),
  1562 => (x"ed",x"49",x"bf",x"ec"),
  1563 => (x"86",x"cc",x"87",x"e6"),
  1564 => (x"bf",x"ec",x"e9",x"c2"),
  1565 => (x"87",x"e5",x"e8",x"49"),
  1566 => (x"c8",x"02",x"9b",x"73"),
  1567 => (x"dc",x"e5",x"c1",x"87"),
  1568 => (x"ca",x"e4",x"c0",x"49"),
  1569 => (x"ec",x"dc",x"ff",x"87"),
  1570 => (x"1e",x"73",x"1e",x"87"),
  1571 => (x"e5",x"c1",x"4b",x"c0"),
  1572 => (x"50",x"c0",x"48",x"c8"),
  1573 => (x"bf",x"ff",x"e6",x"c1"),
  1574 => (x"e6",x"d7",x"ff",x"49"),
  1575 => (x"05",x"98",x"70",x"87"),
  1576 => (x"e2",x"c1",x"87",x"c4"),
  1577 => (x"48",x"73",x"4b",x"ec"),
  1578 => (x"87",x"c9",x"dc",x"ff"),
  1579 => (x"20",x"4d",x"4f",x"52"),
  1580 => (x"64",x"61",x"6f",x"6c"),
  1581 => (x"20",x"67",x"6e",x"69"),
  1582 => (x"6c",x"69",x"61",x"66"),
  1583 => (x"1e",x"00",x"64",x"65"),
  1584 => (x"c1",x"87",x"e3",x"c7"),
  1585 => (x"87",x"c3",x"fe",x"49"),
  1586 => (x"87",x"c3",x"e8",x"fe"),
  1587 => (x"cd",x"02",x"98",x"70"),
  1588 => (x"fe",x"f0",x"fe",x"87"),
  1589 => (x"02",x"98",x"70",x"87"),
  1590 => (x"4a",x"c1",x"87",x"c4"),
  1591 => (x"4a",x"c0",x"87",x"c2"),
  1592 => (x"ce",x"05",x"9a",x"72"),
  1593 => (x"c1",x"1e",x"c0",x"87"),
  1594 => (x"c0",x"49",x"cf",x"e4"),
  1595 => (x"c4",x"87",x"d8",x"ef"),
  1596 => (x"c0",x"87",x"fe",x"86"),
  1597 => (x"da",x"e4",x"c1",x"1e"),
  1598 => (x"ca",x"ef",x"c0",x"49"),
  1599 => (x"fe",x"1e",x"c0",x"87"),
  1600 => (x"49",x"70",x"87",x"c7"),
  1601 => (x"87",x"ff",x"ee",x"c0"),
  1602 => (x"f8",x"87",x"da",x"c3"),
  1603 => (x"53",x"4f",x"26",x"8e"),
  1604 => (x"61",x"66",x"20",x"44"),
  1605 => (x"64",x"65",x"6c",x"69"),
  1606 => (x"6f",x"42",x"00",x"2e"),
  1607 => (x"6e",x"69",x"74",x"6f"),
  1608 => (x"2e",x"2e",x"2e",x"67"),
  1609 => (x"e6",x"c0",x"1e",x"00"),
  1610 => (x"f2",x"c0",x"87",x"e3"),
  1611 => (x"87",x"f6",x"87",x"d3"),
  1612 => (x"c2",x"1e",x"4f",x"26"),
  1613 => (x"c0",x"48",x"c4",x"ea"),
  1614 => (x"ec",x"e9",x"c2",x"78"),
  1615 => (x"fd",x"78",x"c0",x"48"),
  1616 => (x"87",x"e1",x"87",x"fd"),
  1617 => (x"4f",x"26",x"48",x"c0"),
  1618 => (x"00",x"01",x"00",x"00"),
  1619 => (x"20",x"80",x"00",x"00"),
  1620 => (x"74",x"69",x"78",x"45"),
  1621 => (x"42",x"20",x"80",x"00"),
  1622 => (x"00",x"6b",x"63",x"61"),
  1623 => (x"00",x"00",x"10",x"38"),
  1624 => (x"00",x"00",x"2a",x"98"),
  1625 => (x"38",x"00",x"00",x"00"),
  1626 => (x"b6",x"00",x"00",x"10"),
  1627 => (x"00",x"00",x"00",x"2a"),
  1628 => (x"10",x"38",x"00",x"00"),
  1629 => (x"2a",x"d4",x"00",x"00"),
  1630 => (x"00",x"00",x"00",x"00"),
  1631 => (x"00",x"10",x"38",x"00"),
  1632 => (x"00",x"2a",x"f2",x"00"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"00",x"00",x"10",x"38"),
  1635 => (x"00",x"00",x"2b",x"10"),
  1636 => (x"38",x"00",x"00",x"00"),
  1637 => (x"2e",x"00",x"00",x"10"),
  1638 => (x"00",x"00",x"00",x"2b"),
  1639 => (x"10",x"38",x"00",x"00"),
  1640 => (x"2b",x"4c",x"00",x"00"),
  1641 => (x"00",x"00",x"00",x"00"),
  1642 => (x"00",x"12",x"75",x"00"),
  1643 => (x"00",x"00",x"00",x"00"),
  1644 => (x"00",x"00",x"00",x"00"),
  1645 => (x"00",x"00",x"13",x"45"),
  1646 => (x"00",x"00",x"00",x"00"),
  1647 => (x"c3",x"00",x"00",x"00"),
  1648 => (x"53",x"00",x"00",x"19"),
  1649 => (x"49",x"44",x"52",x"4f"),
  1650 => (x"52",x"20",x"54",x"4e"),
  1651 => (x"1e",x"00",x"4d",x"4f"),
  1652 => (x"c0",x"48",x"f0",x"fe"),
  1653 => (x"79",x"09",x"cd",x"78"),
  1654 => (x"1e",x"4f",x"26",x"09"),
  1655 => (x"bf",x"f0",x"fe",x"1e"),
  1656 => (x"26",x"26",x"48",x"7e"),
  1657 => (x"f0",x"fe",x"1e",x"4f"),
  1658 => (x"26",x"78",x"c1",x"48"),
  1659 => (x"f0",x"fe",x"1e",x"4f"),
  1660 => (x"26",x"78",x"c0",x"48"),
  1661 => (x"4a",x"71",x"1e",x"4f"),
  1662 => (x"26",x"52",x"52",x"c0"),
  1663 => (x"5b",x"5e",x"0e",x"4f"),
  1664 => (x"f4",x"0e",x"5d",x"5c"),
  1665 => (x"97",x"4d",x"71",x"86"),
  1666 => (x"a5",x"c1",x"7e",x"6d"),
  1667 => (x"48",x"6c",x"97",x"4c"),
  1668 => (x"6e",x"58",x"a6",x"c8"),
  1669 => (x"a8",x"66",x"c4",x"48"),
  1670 => (x"ff",x"87",x"c5",x"05"),
  1671 => (x"87",x"e6",x"c0",x"48"),
  1672 => (x"c2",x"87",x"ca",x"ff"),
  1673 => (x"6c",x"97",x"49",x"a5"),
  1674 => (x"4b",x"a3",x"71",x"4b"),
  1675 => (x"97",x"4b",x"6b",x"97"),
  1676 => (x"48",x"6e",x"7e",x"6c"),
  1677 => (x"a6",x"c8",x"80",x"c1"),
  1678 => (x"cc",x"98",x"c7",x"58"),
  1679 => (x"97",x"70",x"58",x"a6"),
  1680 => (x"87",x"e1",x"fe",x"7c"),
  1681 => (x"8e",x"f4",x"48",x"73"),
  1682 => (x"4c",x"26",x"4d",x"26"),
  1683 => (x"4f",x"26",x"4b",x"26"),
  1684 => (x"5c",x"5b",x"5e",x"0e"),
  1685 => (x"71",x"86",x"f4",x"0e"),
  1686 => (x"4a",x"66",x"d8",x"4c"),
  1687 => (x"c2",x"9a",x"ff",x"c3"),
  1688 => (x"6c",x"97",x"4b",x"a4"),
  1689 => (x"49",x"a1",x"73",x"49"),
  1690 => (x"6c",x"97",x"51",x"72"),
  1691 => (x"c1",x"48",x"6e",x"7e"),
  1692 => (x"58",x"a6",x"c8",x"80"),
  1693 => (x"a6",x"cc",x"98",x"c7"),
  1694 => (x"f4",x"54",x"70",x"58"),
  1695 => (x"87",x"ca",x"ff",x"8e"),
  1696 => (x"e8",x"fd",x"1e",x"1e"),
  1697 => (x"4a",x"bf",x"e0",x"87"),
  1698 => (x"c0",x"e0",x"c0",x"49"),
  1699 => (x"87",x"cb",x"02",x"99"),
  1700 => (x"ed",x"c2",x"1e",x"72"),
  1701 => (x"f7",x"fe",x"49",x"ea"),
  1702 => (x"fc",x"86",x"c4",x"87"),
  1703 => (x"7e",x"70",x"87",x"fd"),
  1704 => (x"26",x"87",x"c2",x"fd"),
  1705 => (x"c2",x"1e",x"4f",x"26"),
  1706 => (x"fd",x"49",x"ea",x"ed"),
  1707 => (x"ea",x"c1",x"87",x"c7"),
  1708 => (x"da",x"fc",x"49",x"c0"),
  1709 => (x"87",x"f7",x"c3",x"87"),
  1710 => (x"5e",x"0e",x"4f",x"26"),
  1711 => (x"0e",x"5d",x"5c",x"5b"),
  1712 => (x"ed",x"c2",x"4d",x"71"),
  1713 => (x"f4",x"fc",x"49",x"ea"),
  1714 => (x"c0",x"4b",x"70",x"87"),
  1715 => (x"c3",x"04",x"ab",x"b7"),
  1716 => (x"f0",x"c3",x"87",x"c2"),
  1717 => (x"87",x"c9",x"05",x"ab"),
  1718 => (x"48",x"de",x"ee",x"c1"),
  1719 => (x"e3",x"c2",x"78",x"c1"),
  1720 => (x"ab",x"e0",x"c3",x"87"),
  1721 => (x"c1",x"87",x"c9",x"05"),
  1722 => (x"c1",x"48",x"e2",x"ee"),
  1723 => (x"87",x"d4",x"c2",x"78"),
  1724 => (x"bf",x"e2",x"ee",x"c1"),
  1725 => (x"c2",x"87",x"c6",x"02"),
  1726 => (x"c2",x"4c",x"a3",x"c0"),
  1727 => (x"c1",x"4c",x"73",x"87"),
  1728 => (x"02",x"bf",x"de",x"ee"),
  1729 => (x"74",x"87",x"e0",x"c0"),
  1730 => (x"29",x"b7",x"c4",x"49"),
  1731 => (x"fe",x"ef",x"c1",x"91"),
  1732 => (x"cf",x"4a",x"74",x"81"),
  1733 => (x"c1",x"92",x"c2",x"9a"),
  1734 => (x"70",x"30",x"72",x"48"),
  1735 => (x"72",x"ba",x"ff",x"4a"),
  1736 => (x"70",x"98",x"69",x"48"),
  1737 => (x"74",x"87",x"db",x"79"),
  1738 => (x"29",x"b7",x"c4",x"49"),
  1739 => (x"fe",x"ef",x"c1",x"91"),
  1740 => (x"cf",x"4a",x"74",x"81"),
  1741 => (x"c3",x"92",x"c2",x"9a"),
  1742 => (x"70",x"30",x"72",x"48"),
  1743 => (x"b0",x"69",x"48",x"4a"),
  1744 => (x"9d",x"75",x"79",x"70"),
  1745 => (x"87",x"f0",x"c0",x"05"),
  1746 => (x"c8",x"48",x"d0",x"ff"),
  1747 => (x"d4",x"ff",x"78",x"e1"),
  1748 => (x"c1",x"78",x"c5",x"48"),
  1749 => (x"02",x"bf",x"e2",x"ee"),
  1750 => (x"e0",x"c3",x"87",x"c3"),
  1751 => (x"de",x"ee",x"c1",x"78"),
  1752 => (x"87",x"c6",x"02",x"bf"),
  1753 => (x"c3",x"48",x"d4",x"ff"),
  1754 => (x"d4",x"ff",x"78",x"f0"),
  1755 => (x"ff",x"78",x"73",x"48"),
  1756 => (x"e1",x"c8",x"48",x"d0"),
  1757 => (x"78",x"e0",x"c0",x"78"),
  1758 => (x"48",x"e2",x"ee",x"c1"),
  1759 => (x"ee",x"c1",x"78",x"c0"),
  1760 => (x"78",x"c0",x"48",x"de"),
  1761 => (x"49",x"ea",x"ed",x"c2"),
  1762 => (x"70",x"87",x"f2",x"f9"),
  1763 => (x"ab",x"b7",x"c0",x"4b"),
  1764 => (x"87",x"fe",x"fc",x"03"),
  1765 => (x"4d",x"26",x"48",x"c0"),
  1766 => (x"4b",x"26",x"4c",x"26"),
  1767 => (x"00",x"00",x"4f",x"26"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"71",x"1e",x"00",x"00"),
  1770 => (x"cd",x"fc",x"49",x"4a"),
  1771 => (x"1e",x"4f",x"26",x"87"),
  1772 => (x"49",x"72",x"4a",x"c0"),
  1773 => (x"ef",x"c1",x"91",x"c4"),
  1774 => (x"79",x"c0",x"81",x"fe"),
  1775 => (x"b7",x"d0",x"82",x"c1"),
  1776 => (x"87",x"ee",x"04",x"aa"),
  1777 => (x"5e",x"0e",x"4f",x"26"),
  1778 => (x"0e",x"5d",x"5c",x"5b"),
  1779 => (x"dc",x"f8",x"4d",x"71"),
  1780 => (x"c4",x"4a",x"75",x"87"),
  1781 => (x"c1",x"92",x"2a",x"b7"),
  1782 => (x"75",x"82",x"fe",x"ef"),
  1783 => (x"c2",x"9c",x"cf",x"4c"),
  1784 => (x"4b",x"49",x"6a",x"94"),
  1785 => (x"9b",x"c3",x"2b",x"74"),
  1786 => (x"30",x"74",x"48",x"c2"),
  1787 => (x"bc",x"ff",x"4c",x"70"),
  1788 => (x"98",x"71",x"48",x"74"),
  1789 => (x"ec",x"f7",x"7a",x"70"),
  1790 => (x"fe",x"48",x"73",x"87"),
  1791 => (x"00",x"00",x"87",x"d8"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"00",x"00",x"00",x"00"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"00",x"00",x"00",x"00"),
  1806 => (x"00",x"00",x"00",x"00"),
  1807 => (x"ff",x"1e",x"00",x"00"),
  1808 => (x"e1",x"c8",x"48",x"d0"),
  1809 => (x"ff",x"48",x"71",x"78"),
  1810 => (x"26",x"78",x"08",x"d4"),
  1811 => (x"d0",x"ff",x"1e",x"4f"),
  1812 => (x"78",x"e1",x"c8",x"48"),
  1813 => (x"d4",x"ff",x"48",x"71"),
  1814 => (x"66",x"c4",x"78",x"08"),
  1815 => (x"08",x"d4",x"ff",x"48"),
  1816 => (x"1e",x"4f",x"26",x"78"),
  1817 => (x"66",x"c4",x"4a",x"71"),
  1818 => (x"49",x"72",x"1e",x"49"),
  1819 => (x"ff",x"87",x"de",x"ff"),
  1820 => (x"e0",x"c0",x"48",x"d0"),
  1821 => (x"4f",x"26",x"26",x"78"),
  1822 => (x"71",x"1e",x"73",x"1e"),
  1823 => (x"49",x"66",x"c8",x"4b"),
  1824 => (x"c1",x"4a",x"73",x"1e"),
  1825 => (x"ff",x"49",x"a2",x"e0"),
  1826 => (x"c4",x"26",x"87",x"d9"),
  1827 => (x"26",x"4d",x"26",x"87"),
  1828 => (x"26",x"4b",x"26",x"4c"),
  1829 => (x"1e",x"73",x"1e",x"4f"),
  1830 => (x"c2",x"4b",x"4a",x"71"),
  1831 => (x"c8",x"03",x"ab",x"b7"),
  1832 => (x"4a",x"49",x"a3",x"87"),
  1833 => (x"c7",x"9a",x"ff",x"c3"),
  1834 => (x"49",x"a3",x"ce",x"87"),
  1835 => (x"9a",x"ff",x"c3",x"4a"),
  1836 => (x"1e",x"49",x"66",x"c8"),
  1837 => (x"ea",x"fe",x"49",x"72"),
  1838 => (x"d4",x"ff",x"26",x"87"),
  1839 => (x"d4",x"ff",x"1e",x"87"),
  1840 => (x"7a",x"ff",x"c3",x"4a"),
  1841 => (x"c0",x"48",x"d0",x"ff"),
  1842 => (x"7a",x"de",x"78",x"e1"),
  1843 => (x"bf",x"f4",x"ed",x"c2"),
  1844 => (x"c8",x"48",x"49",x"7a"),
  1845 => (x"71",x"7a",x"70",x"28"),
  1846 => (x"70",x"28",x"d0",x"48"),
  1847 => (x"d8",x"48",x"71",x"7a"),
  1848 => (x"ff",x"7a",x"70",x"28"),
  1849 => (x"e0",x"c0",x"48",x"d0"),
  1850 => (x"1e",x"4f",x"26",x"78"),
  1851 => (x"c8",x"48",x"d0",x"ff"),
  1852 => (x"48",x"71",x"78",x"c9"),
  1853 => (x"78",x"08",x"d4",x"ff"),
  1854 => (x"71",x"1e",x"4f",x"26"),
  1855 => (x"87",x"eb",x"49",x"4a"),
  1856 => (x"c8",x"48",x"d0",x"ff"),
  1857 => (x"1e",x"4f",x"26",x"78"),
  1858 => (x"4b",x"71",x"1e",x"73"),
  1859 => (x"bf",x"c4",x"ee",x"c2"),
  1860 => (x"c2",x"87",x"c3",x"02"),
  1861 => (x"d0",x"ff",x"87",x"eb"),
  1862 => (x"78",x"c9",x"c8",x"48"),
  1863 => (x"e0",x"c0",x"49",x"73"),
  1864 => (x"48",x"d4",x"ff",x"b1"),
  1865 => (x"ed",x"c2",x"78",x"71"),
  1866 => (x"78",x"c0",x"48",x"f8"),
  1867 => (x"c5",x"02",x"66",x"c8"),
  1868 => (x"49",x"ff",x"c3",x"87"),
  1869 => (x"49",x"c0",x"87",x"c2"),
  1870 => (x"59",x"c0",x"ee",x"c2"),
  1871 => (x"c6",x"02",x"66",x"cc"),
  1872 => (x"d5",x"d5",x"c5",x"87"),
  1873 => (x"cf",x"87",x"c4",x"4a"),
  1874 => (x"c2",x"4a",x"ff",x"ff"),
  1875 => (x"c2",x"5a",x"c4",x"ee"),
  1876 => (x"c1",x"48",x"c4",x"ee"),
  1877 => (x"26",x"87",x"c4",x"78"),
  1878 => (x"26",x"4c",x"26",x"4d"),
  1879 => (x"0e",x"4f",x"26",x"4b"),
  1880 => (x"5d",x"5c",x"5b",x"5e"),
  1881 => (x"c2",x"4a",x"71",x"0e"),
  1882 => (x"4c",x"bf",x"c0",x"ee"),
  1883 => (x"cb",x"02",x"9a",x"72"),
  1884 => (x"91",x"c8",x"49",x"87"),
  1885 => (x"4b",x"fd",x"f3",x"c1"),
  1886 => (x"87",x"c4",x"83",x"71"),
  1887 => (x"4b",x"fd",x"f7",x"c1"),
  1888 => (x"49",x"13",x"4d",x"c0"),
  1889 => (x"ed",x"c2",x"99",x"74"),
  1890 => (x"ff",x"b9",x"bf",x"fc"),
  1891 => (x"78",x"71",x"48",x"d4"),
  1892 => (x"85",x"2c",x"b7",x"c1"),
  1893 => (x"04",x"ad",x"b7",x"c8"),
  1894 => (x"ed",x"c2",x"87",x"e8"),
  1895 => (x"c8",x"48",x"bf",x"f8"),
  1896 => (x"fc",x"ed",x"c2",x"80"),
  1897 => (x"87",x"ef",x"fe",x"58"),
  1898 => (x"71",x"1e",x"73",x"1e"),
  1899 => (x"9a",x"4a",x"13",x"4b"),
  1900 => (x"72",x"87",x"cb",x"02"),
  1901 => (x"87",x"e7",x"fe",x"49"),
  1902 => (x"05",x"9a",x"4a",x"13"),
  1903 => (x"da",x"fe",x"87",x"f5"),
  1904 => (x"ed",x"c2",x"1e",x"87"),
  1905 => (x"c2",x"49",x"bf",x"f8"),
  1906 => (x"c1",x"48",x"f8",x"ed"),
  1907 => (x"c0",x"c4",x"78",x"a1"),
  1908 => (x"db",x"03",x"a9",x"b7"),
  1909 => (x"48",x"d4",x"ff",x"87"),
  1910 => (x"bf",x"fc",x"ed",x"c2"),
  1911 => (x"f8",x"ed",x"c2",x"78"),
  1912 => (x"ed",x"c2",x"49",x"bf"),
  1913 => (x"a1",x"c1",x"48",x"f8"),
  1914 => (x"b7",x"c0",x"c4",x"78"),
  1915 => (x"87",x"e5",x"04",x"a9"),
  1916 => (x"c8",x"48",x"d0",x"ff"),
  1917 => (x"c4",x"ee",x"c2",x"78"),
  1918 => (x"26",x"78",x"c0",x"48"),
  1919 => (x"00",x"00",x"00",x"4f"),
  1920 => (x"00",x"00",x"00",x"00"),
  1921 => (x"00",x"00",x"00",x"00"),
  1922 => (x"00",x"00",x"5f",x"5f"),
  1923 => (x"03",x"03",x"00",x"00"),
  1924 => (x"00",x"03",x"03",x"00"),
  1925 => (x"7f",x"7f",x"14",x"00"),
  1926 => (x"14",x"7f",x"7f",x"14"),
  1927 => (x"2e",x"24",x"00",x"00"),
  1928 => (x"12",x"3a",x"6b",x"6b"),
  1929 => (x"36",x"6a",x"4c",x"00"),
  1930 => (x"32",x"56",x"6c",x"18"),
  1931 => (x"4f",x"7e",x"30",x"00"),
  1932 => (x"68",x"3a",x"77",x"59"),
  1933 => (x"04",x"00",x"00",x"40"),
  1934 => (x"00",x"00",x"03",x"07"),
  1935 => (x"1c",x"00",x"00",x"00"),
  1936 => (x"00",x"41",x"63",x"3e"),
  1937 => (x"41",x"00",x"00",x"00"),
  1938 => (x"00",x"1c",x"3e",x"63"),
  1939 => (x"3e",x"2a",x"08",x"00"),
  1940 => (x"2a",x"3e",x"1c",x"1c"),
  1941 => (x"08",x"08",x"00",x"08"),
  1942 => (x"08",x"08",x"3e",x"3e"),
  1943 => (x"80",x"00",x"00",x"00"),
  1944 => (x"00",x"00",x"60",x"e0"),
  1945 => (x"08",x"08",x"00",x"00"),
  1946 => (x"08",x"08",x"08",x"08"),
  1947 => (x"00",x"00",x"00",x"00"),
  1948 => (x"00",x"00",x"60",x"60"),
  1949 => (x"30",x"60",x"40",x"00"),
  1950 => (x"03",x"06",x"0c",x"18"),
  1951 => (x"7f",x"3e",x"00",x"01"),
  1952 => (x"3e",x"7f",x"4d",x"59"),
  1953 => (x"06",x"04",x"00",x"00"),
  1954 => (x"00",x"00",x"7f",x"7f"),
  1955 => (x"63",x"42",x"00",x"00"),
  1956 => (x"46",x"4f",x"59",x"71"),
  1957 => (x"63",x"22",x"00",x"00"),
  1958 => (x"36",x"7f",x"49",x"49"),
  1959 => (x"16",x"1c",x"18",x"00"),
  1960 => (x"10",x"7f",x"7f",x"13"),
  1961 => (x"67",x"27",x"00",x"00"),
  1962 => (x"39",x"7d",x"45",x"45"),
  1963 => (x"7e",x"3c",x"00",x"00"),
  1964 => (x"30",x"79",x"49",x"4b"),
  1965 => (x"01",x"01",x"00",x"00"),
  1966 => (x"07",x"0f",x"79",x"71"),
  1967 => (x"7f",x"36",x"00",x"00"),
  1968 => (x"36",x"7f",x"49",x"49"),
  1969 => (x"4f",x"06",x"00",x"00"),
  1970 => (x"1e",x"3f",x"69",x"49"),
  1971 => (x"00",x"00",x"00",x"00"),
  1972 => (x"00",x"00",x"66",x"66"),
  1973 => (x"80",x"00",x"00",x"00"),
  1974 => (x"00",x"00",x"66",x"e6"),
  1975 => (x"08",x"08",x"00",x"00"),
  1976 => (x"22",x"22",x"14",x"14"),
  1977 => (x"14",x"14",x"00",x"00"),
  1978 => (x"14",x"14",x"14",x"14"),
  1979 => (x"22",x"22",x"00",x"00"),
  1980 => (x"08",x"08",x"14",x"14"),
  1981 => (x"03",x"02",x"00",x"00"),
  1982 => (x"06",x"0f",x"59",x"51"),
  1983 => (x"41",x"7f",x"3e",x"00"),
  1984 => (x"1e",x"1f",x"55",x"5d"),
  1985 => (x"7f",x"7e",x"00",x"00"),
  1986 => (x"7e",x"7f",x"09",x"09"),
  1987 => (x"7f",x"7f",x"00",x"00"),
  1988 => (x"36",x"7f",x"49",x"49"),
  1989 => (x"3e",x"1c",x"00",x"00"),
  1990 => (x"41",x"41",x"41",x"63"),
  1991 => (x"7f",x"7f",x"00",x"00"),
  1992 => (x"1c",x"3e",x"63",x"41"),
  1993 => (x"7f",x"7f",x"00",x"00"),
  1994 => (x"41",x"41",x"49",x"49"),
  1995 => (x"7f",x"7f",x"00",x"00"),
  1996 => (x"01",x"01",x"09",x"09"),
  1997 => (x"7f",x"3e",x"00",x"00"),
  1998 => (x"7a",x"7b",x"49",x"41"),
  1999 => (x"7f",x"7f",x"00",x"00"),
  2000 => (x"7f",x"7f",x"08",x"08"),
  2001 => (x"41",x"00",x"00",x"00"),
  2002 => (x"00",x"41",x"7f",x"7f"),
  2003 => (x"60",x"20",x"00",x"00"),
  2004 => (x"3f",x"7f",x"40",x"40"),
  2005 => (x"08",x"7f",x"7f",x"00"),
  2006 => (x"41",x"63",x"36",x"1c"),
  2007 => (x"7f",x"7f",x"00",x"00"),
  2008 => (x"40",x"40",x"40",x"40"),
  2009 => (x"06",x"7f",x"7f",x"00"),
  2010 => (x"7f",x"7f",x"06",x"0c"),
  2011 => (x"06",x"7f",x"7f",x"00"),
  2012 => (x"7f",x"7f",x"18",x"0c"),
  2013 => (x"7f",x"3e",x"00",x"00"),
  2014 => (x"3e",x"7f",x"41",x"41"),
  2015 => (x"7f",x"7f",x"00",x"00"),
  2016 => (x"06",x"0f",x"09",x"09"),
  2017 => (x"41",x"7f",x"3e",x"00"),
  2018 => (x"40",x"7e",x"7f",x"61"),
  2019 => (x"7f",x"7f",x"00",x"00"),
  2020 => (x"66",x"7f",x"19",x"09"),
  2021 => (x"6f",x"26",x"00",x"00"),
  2022 => (x"32",x"7b",x"59",x"4d"),
  2023 => (x"01",x"01",x"00",x"00"),
  2024 => (x"01",x"01",x"7f",x"7f"),
  2025 => (x"7f",x"3f",x"00",x"00"),
  2026 => (x"3f",x"7f",x"40",x"40"),
  2027 => (x"3f",x"0f",x"00",x"00"),
  2028 => (x"0f",x"3f",x"70",x"70"),
  2029 => (x"30",x"7f",x"7f",x"00"),
  2030 => (x"7f",x"7f",x"30",x"18"),
  2031 => (x"36",x"63",x"41",x"00"),
  2032 => (x"63",x"36",x"1c",x"1c"),
  2033 => (x"06",x"03",x"01",x"41"),
  2034 => (x"03",x"06",x"7c",x"7c"),
  2035 => (x"59",x"71",x"61",x"01"),
  2036 => (x"41",x"43",x"47",x"4d"),
  2037 => (x"7f",x"00",x"00",x"00"),
  2038 => (x"00",x"41",x"41",x"7f"),
  2039 => (x"06",x"03",x"01",x"00"),
  2040 => (x"60",x"30",x"18",x"0c"),
  2041 => (x"41",x"00",x"00",x"40"),
  2042 => (x"00",x"7f",x"7f",x"41"),
  2043 => (x"06",x"0c",x"08",x"00"),
  2044 => (x"08",x"0c",x"06",x"03"),
  2045 => (x"80",x"80",x"80",x"00"),
  2046 => (x"80",x"80",x"80",x"80"),
  2047 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

