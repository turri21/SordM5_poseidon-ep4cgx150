library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c8efc287",
    12 => x"86c0c84e",
    13 => x"49c8efc2",
    14 => x"48d4dcc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e7e3",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34972",
    82 => x"c27c7199",
    83 => x"05bfd4dc",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"c329d849",
    88 => x"7c7199ff",
    89 => x"d04966d0",
    90 => x"99ffc329",
    91 => x"66d07c71",
    92 => x"c329c849",
    93 => x"7c7199ff",
    94 => x"c34966d0",
    95 => x"7c7199ff",
    96 => x"29d04972",
    97 => x"7199ffc3",
    98 => x"c94b6c7c",
    99 => x"c34dfff0",
   100 => x"d005abff",
   101 => x"7cffc387",
   102 => x"8dc14b6c",
   103 => x"c387c602",
   104 => x"f002abff",
   105 => x"fe487387",
   106 => x"c01e87c7",
   107 => x"48d4ff49",
   108 => x"c178ffc3",
   109 => x"b7c8c381",
   110 => x"87f104a9",
   111 => x"731e4f26",
   112 => x"c487e71e",
   113 => x"c04bdff8",
   114 => x"f0ffc01e",
   115 => x"fd49f7c1",
   116 => x"86c487e7",
   117 => x"c005a8c1",
   118 => x"d4ff87ea",
   119 => x"78ffc348",
   120 => x"c0c0c0c1",
   121 => x"c01ec0c0",
   122 => x"e9c1f0e1",
   123 => x"87c9fd49",
   124 => x"987086c4",
   125 => x"ff87ca05",
   126 => x"ffc348d4",
   127 => x"cb48c178",
   128 => x"87e6fe87",
   129 => x"fe058bc1",
   130 => x"48c087fd",
   131 => x"1e87e6fc",
   132 => x"d4ff1e73",
   133 => x"78ffc348",
   134 => x"1ec04bd3",
   135 => x"c1f0ffc0",
   136 => x"d4fc49c1",
   137 => x"7086c487",
   138 => x"87ca0598",
   139 => x"c348d4ff",
   140 => x"48c178ff",
   141 => x"f1fd87cb",
   142 => x"058bc187",
   143 => x"c087dbff",
   144 => x"87f1fb48",
   145 => x"5c5b5e0e",
   146 => x"4cd4ff0e",
   147 => x"c687dbfd",
   148 => x"e1c01eea",
   149 => x"49c8c1f0",
   150 => x"c487defb",
   151 => x"02a8c186",
   152 => x"eafe87c8",
   153 => x"c148c087",
   154 => x"dafa87e2",
   155 => x"cf497087",
   156 => x"c699ffff",
   157 => x"c802a9ea",
   158 => x"87d3fe87",
   159 => x"cbc148c0",
   160 => x"7cffc387",
   161 => x"fc4bf1c0",
   162 => x"987087f4",
   163 => x"87ebc002",
   164 => x"ffc01ec0",
   165 => x"49fac1f0",
   166 => x"c487defa",
   167 => x"05987086",
   168 => x"ffc387d9",
   169 => x"c3496c7c",
   170 => x"7c7c7cff",
   171 => x"99c0c17c",
   172 => x"c187c402",
   173 => x"c087d548",
   174 => x"c287d148",
   175 => x"87c405ab",
   176 => x"87c848c0",
   177 => x"fe058bc1",
   178 => x"48c087fd",
   179 => x"1e87e4f9",
   180 => x"dcc21e73",
   181 => x"78c148d4",
   182 => x"d0ff4bc7",
   183 => x"fb78c248",
   184 => x"d0ff87c8",
   185 => x"c078c348",
   186 => x"d0e5c01e",
   187 => x"f949c0c1",
   188 => x"86c487c7",
   189 => x"c105a8c1",
   190 => x"abc24b87",
   191 => x"c087c505",
   192 => x"87f9c048",
   193 => x"ff058bc1",
   194 => x"f7fc87d0",
   195 => x"d8dcc287",
   196 => x"05987058",
   197 => x"1ec187cd",
   198 => x"c1f0ffc0",
   199 => x"d8f849d0",
   200 => x"ff86c487",
   201 => x"ffc348d4",
   202 => x"87dec478",
   203 => x"58dcdcc2",
   204 => x"c248d0ff",
   205 => x"48d4ff78",
   206 => x"c178ffc3",
   207 => x"87f5f748",
   208 => x"5c5b5e0e",
   209 => x"4a710e5d",
   210 => x"ff4dffc3",
   211 => x"7c754cd4",
   212 => x"c448d0ff",
   213 => x"7c7578c3",
   214 => x"ffc01e72",
   215 => x"49d8c1f0",
   216 => x"c487d6f7",
   217 => x"02987086",
   218 => x"48c187c5",
   219 => x"7587f0c0",
   220 => x"7cfec37c",
   221 => x"d41ec0c8",
   222 => x"faf44966",
   223 => x"7586c487",
   224 => x"757c757c",
   225 => x"e0dad87c",
   226 => x"6c7c754b",
   227 => x"c5059949",
   228 => x"058bc187",
   229 => x"7c7587f3",
   230 => x"c248d0ff",
   231 => x"f648c078",
   232 => x"5e0e87cf",
   233 => x"0e5d5c5b",
   234 => x"4cc04b71",
   235 => x"dfcdeec5",
   236 => x"48d4ff4a",
   237 => x"6878ffc3",
   238 => x"a9fec349",
   239 => x"87fdc005",
   240 => x"9b734d70",
   241 => x"d087cc02",
   242 => x"49731e66",
   243 => x"c487cff4",
   244 => x"ff87d686",
   245 => x"d1c448d0",
   246 => x"7dffc378",
   247 => x"c14866d0",
   248 => x"58a6d488",
   249 => x"f0059870",
   250 => x"48d4ff87",
   251 => x"7878ffc3",
   252 => x"c5059b73",
   253 => x"48d0ff87",
   254 => x"4ac178d0",
   255 => x"058ac14c",
   256 => x"7487eefe",
   257 => x"87e9f448",
   258 => x"711e731e",
   259 => x"ff4bc04a",
   260 => x"ffc348d4",
   261 => x"48d0ff78",
   262 => x"ff78c3c4",
   263 => x"ffc348d4",
   264 => x"c01e7278",
   265 => x"d1c1f0ff",
   266 => x"87cdf449",
   267 => x"987086c4",
   268 => x"c887d205",
   269 => x"66cc1ec0",
   270 => x"87e6fd49",
   271 => x"4b7086c4",
   272 => x"c248d0ff",
   273 => x"f3487378",
   274 => x"5e0e87eb",
   275 => x"0e5d5c5b",
   276 => x"ffc01ec0",
   277 => x"49c9c1f0",
   278 => x"d287def3",
   279 => x"dcdcc21e",
   280 => x"87fefc49",
   281 => x"4cc086c8",
   282 => x"b7d284c1",
   283 => x"87f804ac",
   284 => x"97dcdcc2",
   285 => x"c0c349bf",
   286 => x"a9c0c199",
   287 => x"87e7c005",
   288 => x"97e3dcc2",
   289 => x"31d049bf",
   290 => x"97e4dcc2",
   291 => x"32c84abf",
   292 => x"dcc2b172",
   293 => x"4abf97e5",
   294 => x"cf4c71b1",
   295 => x"9cffffff",
   296 => x"34ca84c1",
   297 => x"c287e7c1",
   298 => x"bf97e5dc",
   299 => x"c631c149",
   300 => x"e6dcc299",
   301 => x"c74abf97",
   302 => x"b1722ab7",
   303 => x"97e1dcc2",
   304 => x"cf4d4abf",
   305 => x"e2dcc29d",
   306 => x"c34abf97",
   307 => x"c232ca9a",
   308 => x"bf97e3dc",
   309 => x"7333c24b",
   310 => x"e4dcc2b2",
   311 => x"c34bbf97",
   312 => x"b7c69bc0",
   313 => x"c2b2732b",
   314 => x"7148c181",
   315 => x"c1497030",
   316 => x"70307548",
   317 => x"c14c724d",
   318 => x"c8947184",
   319 => x"06adb7c0",
   320 => x"34c187cc",
   321 => x"c0c82db7",
   322 => x"ff01adb7",
   323 => x"487487f4",
   324 => x"0e87def0",
   325 => x"5d5c5b5e",
   326 => x"c286f80e",
   327 => x"c048c2e5",
   328 => x"fadcc278",
   329 => x"fb49c01e",
   330 => x"86c487de",
   331 => x"c5059870",
   332 => x"c948c087",
   333 => x"4dc087ce",
   334 => x"f2c07ec1",
   335 => x"c249bfed",
   336 => x"714af0dd",
   337 => x"e0ec4bc8",
   338 => x"05987087",
   339 => x"7ec087c2",
   340 => x"bfe9f2c0",
   341 => x"ccdec249",
   342 => x"4bc8714a",
   343 => x"7087caec",
   344 => x"87c20598",
   345 => x"026e7ec0",
   346 => x"c287fdc0",
   347 => x"4dbfc0e4",
   348 => x"9ff8e4c2",
   349 => x"c5487ebf",
   350 => x"05a8ead6",
   351 => x"e4c287c7",
   352 => x"ce4dbfc0",
   353 => x"ca486e87",
   354 => x"02a8d5e9",
   355 => x"48c087c5",
   356 => x"c287f1c7",
   357 => x"751efadc",
   358 => x"87ecf949",
   359 => x"987086c4",
   360 => x"c087c505",
   361 => x"87dcc748",
   362 => x"bfe9f2c0",
   363 => x"ccdec249",
   364 => x"4bc8714a",
   365 => x"7087f2ea",
   366 => x"87c80598",
   367 => x"48c2e5c2",
   368 => x"87da78c1",
   369 => x"bfedf2c0",
   370 => x"f0ddc249",
   371 => x"4bc8714a",
   372 => x"7087d6ea",
   373 => x"c5c00298",
   374 => x"c648c087",
   375 => x"e4c287e6",
   376 => x"49bf97f8",
   377 => x"05a9d5c1",
   378 => x"c287cdc0",
   379 => x"bf97f9e4",
   380 => x"a9eac249",
   381 => x"87c5c002",
   382 => x"c7c648c0",
   383 => x"fadcc287",
   384 => x"487ebf97",
   385 => x"02a8e9c3",
   386 => x"6e87cec0",
   387 => x"a8ebc348",
   388 => x"87c5c002",
   389 => x"ebc548c0",
   390 => x"c5ddc287",
   391 => x"9949bf97",
   392 => x"87ccc005",
   393 => x"97c6ddc2",
   394 => x"a9c249bf",
   395 => x"87c5c002",
   396 => x"cfc548c0",
   397 => x"c7ddc287",
   398 => x"c248bf97",
   399 => x"7058fee4",
   400 => x"88c1484c",
   401 => x"58c2e5c2",
   402 => x"97c8ddc2",
   403 => x"817549bf",
   404 => x"97c9ddc2",
   405 => x"32c84abf",
   406 => x"c27ea172",
   407 => x"6e48cfe9",
   408 => x"caddc278",
   409 => x"c848bf97",
   410 => x"e5c258a6",
   411 => x"c202bfc2",
   412 => x"f2c087d4",
   413 => x"c249bfe9",
   414 => x"714accde",
   415 => x"e8e74bc8",
   416 => x"02987087",
   417 => x"c087c5c0",
   418 => x"87f8c348",
   419 => x"bffae4c2",
   420 => x"e3e9c24c",
   421 => x"dfddc25c",
   422 => x"c849bf97",
   423 => x"deddc231",
   424 => x"a14abf97",
   425 => x"e0ddc249",
   426 => x"d04abf97",
   427 => x"49a17232",
   428 => x"97e1ddc2",
   429 => x"32d84abf",
   430 => x"c449a172",
   431 => x"e9c29166",
   432 => x"c281bfcf",
   433 => x"c259d7e9",
   434 => x"bf97e7dd",
   435 => x"c232c84a",
   436 => x"bf97e6dd",
   437 => x"c24aa24b",
   438 => x"bf97e8dd",
   439 => x"7333d04b",
   440 => x"ddc24aa2",
   441 => x"4bbf97e9",
   442 => x"33d89bcf",
   443 => x"c24aa273",
   444 => x"c25adbe9",
   445 => x"4abfd7e9",
   446 => x"92748ac2",
   447 => x"48dbe9c2",
   448 => x"c178a172",
   449 => x"ddc287ca",
   450 => x"49bf97cc",
   451 => x"ddc231c8",
   452 => x"4abf97cb",
   453 => x"e5c249a1",
   454 => x"e5c259ca",
   455 => x"c549bfc6",
   456 => x"81ffc731",
   457 => x"e9c229c9",
   458 => x"ddc259e3",
   459 => x"4abf97d1",
   460 => x"ddc232c8",
   461 => x"4bbf97d0",
   462 => x"66c44aa2",
   463 => x"c2826e92",
   464 => x"c25adfe9",
   465 => x"c048d7e9",
   466 => x"d3e9c278",
   467 => x"78a17248",
   468 => x"48e3e9c2",
   469 => x"bfd7e9c2",
   470 => x"e7e9c278",
   471 => x"dbe9c248",
   472 => x"e5c278bf",
   473 => x"c002bfc2",
   474 => x"487487c9",
   475 => x"7e7030c4",
   476 => x"c287c9c0",
   477 => x"48bfdfe9",
   478 => x"7e7030c4",
   479 => x"48c6e5c2",
   480 => x"48c1786e",
   481 => x"4d268ef8",
   482 => x"4b264c26",
   483 => x"5e0e4f26",
   484 => x"0e5d5c5b",
   485 => x"e5c24a71",
   486 => x"cb02bfc2",
   487 => x"c74b7287",
   488 => x"c14c722b",
   489 => x"87c99cff",
   490 => x"2bc84b72",
   491 => x"ffc34c72",
   492 => x"cfe9c29c",
   493 => x"f2c083bf",
   494 => x"02abbfe5",
   495 => x"f2c087d9",
   496 => x"dcc25be9",
   497 => x"49731efa",
   498 => x"c487fdf0",
   499 => x"05987086",
   500 => x"48c087c5",
   501 => x"c287e6c0",
   502 => x"02bfc2e5",
   503 => x"497487d2",
   504 => x"dcc291c4",
   505 => x"4d6981fa",
   506 => x"ffffffcf",
   507 => x"87cb9dff",
   508 => x"91c24974",
   509 => x"81fadcc2",
   510 => x"754d699f",
   511 => x"87c6fe48",
   512 => x"5c5b5e0e",
   513 => x"86f80e5d",
   514 => x"059c4c71",
   515 => x"48c087c5",
   516 => x"c887c2c3",
   517 => x"486e7ea4",
   518 => x"66d878c0",
   519 => x"d887c702",
   520 => x"05bf9766",
   521 => x"48c087c5",
   522 => x"c087eac2",
   523 => x"4949c11e",
   524 => x"c487d7ca",
   525 => x"9d4d7086",
   526 => x"87c2c102",
   527 => x"4acae5c2",
   528 => x"e04966d8",
   529 => x"987087c8",
   530 => x"87f2c002",
   531 => x"66d84a75",
   532 => x"e04bcb49",
   533 => x"987087ed",
   534 => x"87e2c002",
   535 => x"9d751ec0",
   536 => x"c887c702",
   537 => x"78c048a6",
   538 => x"a6c887c5",
   539 => x"c878c148",
   540 => x"d5c94966",
   541 => x"7086c487",
   542 => x"fe059d4d",
   543 => x"9d7587fe",
   544 => x"87cfc102",
   545 => x"6e49a5dc",
   546 => x"da786948",
   547 => x"a6c449a5",
   548 => x"78a4c448",
   549 => x"c448699f",
   550 => x"c2780866",
   551 => x"02bfc2e5",
   552 => x"a5d487d2",
   553 => x"49699f49",
   554 => x"99ffffc0",
   555 => x"30d04871",
   556 => x"87c27e70",
   557 => x"496e7ec0",
   558 => x"bf66c448",
   559 => x"0866c480",
   560 => x"cc7cc078",
   561 => x"66c449a4",
   562 => x"a4d079bf",
   563 => x"c179c049",
   564 => x"c087c248",
   565 => x"fa8ef848",
   566 => x"5e0e87ec",
   567 => x"0e5d5c5b",
   568 => x"029c4c71",
   569 => x"c887cac1",
   570 => x"026949a4",
   571 => x"d087c2c1",
   572 => x"496c4a66",
   573 => x"5aa6d482",
   574 => x"b94d66d0",
   575 => x"bffee4c2",
   576 => x"72baff4a",
   577 => x"02997199",
   578 => x"c487e4c0",
   579 => x"496b4ba4",
   580 => x"7087fbf9",
   581 => x"fae4c27b",
   582 => x"816c49bf",
   583 => x"b9757c71",
   584 => x"bffee4c2",
   585 => x"72baff4a",
   586 => x"05997199",
   587 => x"7587dcff",
   588 => x"87d2f97c",
   589 => x"711e731e",
   590 => x"c7029b4b",
   591 => x"49a3c887",
   592 => x"87c50569",
   593 => x"f7c048c0",
   594 => x"d3e9c287",
   595 => x"a3c44abf",
   596 => x"c2496949",
   597 => x"fae4c289",
   598 => x"a27191bf",
   599 => x"fee4c24a",
   600 => x"996b49bf",
   601 => x"c04aa271",
   602 => x"c85ae9f2",
   603 => x"49721e66",
   604 => x"c487d5ea",
   605 => x"05987086",
   606 => x"48c087c4",
   607 => x"48c187c2",
   608 => x"1e87c7f8",
   609 => x"4b711e73",
   610 => x"87c7029b",
   611 => x"6949a3c8",
   612 => x"c087c505",
   613 => x"87f7c048",
   614 => x"bfd3e9c2",
   615 => x"49a3c44a",
   616 => x"89c24969",
   617 => x"bffae4c2",
   618 => x"4aa27191",
   619 => x"bffee4c2",
   620 => x"71996b49",
   621 => x"f2c04aa2",
   622 => x"66c85ae9",
   623 => x"e549721e",
   624 => x"86c487fe",
   625 => x"c4059870",
   626 => x"c248c087",
   627 => x"f648c187",
   628 => x"5e0e87f8",
   629 => x"0e5d5c5b",
   630 => x"d44b711e",
   631 => x"9b734d66",
   632 => x"87ccc102",
   633 => x"6949a3c8",
   634 => x"87c4c102",
   635 => x"c24ca3d0",
   636 => x"49bffee4",
   637 => x"4a6cb9ff",
   638 => x"66d47e99",
   639 => x"87cd06a9",
   640 => x"cc7c7bc0",
   641 => x"a3c44aa3",
   642 => x"ca796a49",
   643 => x"f8497287",
   644 => x"66d499c0",
   645 => x"758d714d",
   646 => x"7129c949",
   647 => x"fa49731e",
   648 => x"dcc287f8",
   649 => x"49731efa",
   650 => x"c887c9fc",
   651 => x"7c66d486",
   652 => x"87d2f526",
   653 => x"711e731e",
   654 => x"c0029b4b",
   655 => x"e9c287e4",
   656 => x"4a735be7",
   657 => x"e4c28ac2",
   658 => x"9249bffa",
   659 => x"bfd3e9c2",
   660 => x"c2807248",
   661 => x"7158ebe9",
   662 => x"c230c448",
   663 => x"c058cae5",
   664 => x"e9c287ed",
   665 => x"e9c248e3",
   666 => x"c278bfd7",
   667 => x"c248e7e9",
   668 => x"78bfdbe9",
   669 => x"bfc2e5c2",
   670 => x"c287c902",
   671 => x"49bffae4",
   672 => x"87c731c4",
   673 => x"bfdfe9c2",
   674 => x"c231c449",
   675 => x"f359cae5",
   676 => x"5e0e87f8",
   677 => x"710e5c5b",
   678 => x"724bc04a",
   679 => x"e1c0029a",
   680 => x"49a2da87",
   681 => x"c24b699f",
   682 => x"02bfc2e5",
   683 => x"a2d487cf",
   684 => x"49699f49",
   685 => x"ffffc04c",
   686 => x"c234d09c",
   687 => x"744cc087",
   688 => x"4973b349",
   689 => x"f287edfd",
   690 => x"5e0e87fe",
   691 => x"0e5d5c5b",
   692 => x"4a7186f4",
   693 => x"9a727ec0",
   694 => x"c287d802",
   695 => x"c048f6dc",
   696 => x"eedcc278",
   697 => x"e7e9c248",
   698 => x"dcc278bf",
   699 => x"e9c248f2",
   700 => x"c278bfe3",
   701 => x"c048d7e5",
   702 => x"c6e5c250",
   703 => x"dcc249bf",
   704 => x"714abff6",
   705 => x"c9c403aa",
   706 => x"cf497287",
   707 => x"e9c00599",
   708 => x"e5f2c087",
   709 => x"eedcc248",
   710 => x"dcc278bf",
   711 => x"dcc21efa",
   712 => x"c249bfee",
   713 => x"c148eedc",
   714 => x"e37178a1",
   715 => x"86c487da",
   716 => x"48e1f2c0",
   717 => x"78fadcc2",
   718 => x"f2c087cc",
   719 => x"c048bfe1",
   720 => x"f2c080e0",
   721 => x"dcc258e5",
   722 => x"c148bff6",
   723 => x"fadcc280",
   724 => x"0ca12758",
   725 => x"97bf0000",
   726 => x"029d4dbf",
   727 => x"c387e3c2",
   728 => x"c202ade5",
   729 => x"f2c087dc",
   730 => x"cb4bbfe1",
   731 => x"4c1149a3",
   732 => x"c105accf",
   733 => x"497587d2",
   734 => x"89c199df",
   735 => x"e5c291cd",
   736 => x"a3c181ca",
   737 => x"c351124a",
   738 => x"51124aa3",
   739 => x"124aa3c5",
   740 => x"4aa3c751",
   741 => x"a3c95112",
   742 => x"ce51124a",
   743 => x"51124aa3",
   744 => x"124aa3d0",
   745 => x"4aa3d251",
   746 => x"a3d45112",
   747 => x"d651124a",
   748 => x"51124aa3",
   749 => x"124aa3d8",
   750 => x"4aa3dc51",
   751 => x"a3de5112",
   752 => x"c151124a",
   753 => x"87fac07e",
   754 => x"99c84974",
   755 => x"87ebc005",
   756 => x"99d04974",
   757 => x"dc87d105",
   758 => x"cbc00266",
   759 => x"dc497387",
   760 => x"98700f66",
   761 => x"87d3c002",
   762 => x"c6c0056e",
   763 => x"cae5c287",
   764 => x"c050c048",
   765 => x"48bfe1f2",
   766 => x"c287e1c2",
   767 => x"c048d7e5",
   768 => x"e5c27e50",
   769 => x"c249bfc6",
   770 => x"4abff6dc",
   771 => x"fb04aa71",
   772 => x"e9c287f7",
   773 => x"c005bfe7",
   774 => x"e5c287c8",
   775 => x"c102bfc2",
   776 => x"dcc287f8",
   777 => x"ed49bff2",
   778 => x"497087e4",
   779 => x"59f6dcc2",
   780 => x"c248a6c4",
   781 => x"78bff2dc",
   782 => x"bfc2e5c2",
   783 => x"87d8c002",
   784 => x"cf4966c4",
   785 => x"f8ffffff",
   786 => x"c002a999",
   787 => x"4cc087c5",
   788 => x"c187e1c0",
   789 => x"87dcc04c",
   790 => x"cf4966c4",
   791 => x"a999f8ff",
   792 => x"87c8c002",
   793 => x"c048a6c8",
   794 => x"87c5c078",
   795 => x"c148a6c8",
   796 => x"4c66c878",
   797 => x"c0059c74",
   798 => x"66c487e0",
   799 => x"c289c249",
   800 => x"4abffae4",
   801 => x"d3e9c291",
   802 => x"dcc24abf",
   803 => x"a17248ee",
   804 => x"f6dcc278",
   805 => x"f978c048",
   806 => x"48c087df",
   807 => x"e5eb8ef4",
   808 => x"00000087",
   809 => x"ffffff00",
   810 => x"000cb1ff",
   811 => x"000cba00",
   812 => x"54414600",
   813 => x"20203233",
   814 => x"41460020",
   815 => x"20363154",
   816 => x"1e002020",
   817 => x"c348d4ff",
   818 => x"486878ff",
   819 => x"ff1e4f26",
   820 => x"ffc348d4",
   821 => x"48d0ff78",
   822 => x"ff78e1c0",
   823 => x"78d448d4",
   824 => x"48ebe9c2",
   825 => x"50bfd4ff",
   826 => x"ff1e4f26",
   827 => x"e0c048d0",
   828 => x"1e4f2678",
   829 => x"7087ccff",
   830 => x"c6029949",
   831 => x"a9fbc087",
   832 => x"7187f105",
   833 => x"0e4f2648",
   834 => x"0e5c5b5e",
   835 => x"4cc04b71",
   836 => x"7087f0fe",
   837 => x"c0029949",
   838 => x"ecc087f9",
   839 => x"f2c002a9",
   840 => x"a9fbc087",
   841 => x"87ebc002",
   842 => x"acb766cc",
   843 => x"d087c703",
   844 => x"87c20266",
   845 => x"99715371",
   846 => x"c187c202",
   847 => x"87c3fe84",
   848 => x"02994970",
   849 => x"ecc087cd",
   850 => x"87c702a9",
   851 => x"05a9fbc0",
   852 => x"d087d5ff",
   853 => x"87c30266",
   854 => x"c07b97c0",
   855 => x"c405a9ec",
   856 => x"c54a7487",
   857 => x"c04a7487",
   858 => x"48728a0a",
   859 => x"4d2687c2",
   860 => x"4b264c26",
   861 => x"fd1e4f26",
   862 => x"497087c9",
   863 => x"aaf0c04a",
   864 => x"c087c904",
   865 => x"c301aaf9",
   866 => x"8af0c087",
   867 => x"04aac1c1",
   868 => x"dac187c9",
   869 => x"87c301aa",
   870 => x"728af7c0",
   871 => x"0e4f2648",
   872 => x"0e5c5b5e",
   873 => x"d4ff4a71",
   874 => x"c049724b",
   875 => x"4c7087e7",
   876 => x"87c2029c",
   877 => x"d0ff8cc1",
   878 => x"c178c548",
   879 => x"49747bd5",
   880 => x"e5c131c6",
   881 => x"4abf97c8",
   882 => x"70b07148",
   883 => x"48d0ff7b",
   884 => x"dbfe78c4",
   885 => x"5b5e0e87",
   886 => x"f80e5d5c",
   887 => x"c04c7186",
   888 => x"87eafb7e",
   889 => x"fac04bc0",
   890 => x"49bf97c2",
   891 => x"cf04a9c0",
   892 => x"87fffb87",
   893 => x"fac083c1",
   894 => x"49bf97c2",
   895 => x"87f106ab",
   896 => x"97c2fac0",
   897 => x"87cf02bf",
   898 => x"7087f8fa",
   899 => x"c6029949",
   900 => x"a9ecc087",
   901 => x"c087f105",
   902 => x"87e7fa4b",
   903 => x"e2fa4d70",
   904 => x"58a6c887",
   905 => x"7087dcfa",
   906 => x"c883c14a",
   907 => x"699749a4",
   908 => x"c702ad49",
   909 => x"adffc087",
   910 => x"87e7c005",
   911 => x"9749a4c9",
   912 => x"66c44969",
   913 => x"87c702a9",
   914 => x"a8ffc048",
   915 => x"ca87d405",
   916 => x"699749a4",
   917 => x"c602aa49",
   918 => x"aaffc087",
   919 => x"c187c405",
   920 => x"c087d07e",
   921 => x"c602adec",
   922 => x"adfbc087",
   923 => x"c087c405",
   924 => x"6e7ec14b",
   925 => x"87e1fe02",
   926 => x"7387eff9",
   927 => x"fb8ef848",
   928 => x"0e0087ec",
   929 => x"5d5c5b5e",
   930 => x"7186f80e",
   931 => x"4bd4ff4d",
   932 => x"e9c21e75",
   933 => x"e7e549f0",
   934 => x"7086c487",
   935 => x"ccc40298",
   936 => x"48a6c487",
   937 => x"bfcae5c1",
   938 => x"fb497578",
   939 => x"d0ff87f1",
   940 => x"c178c548",
   941 => x"4ac07bd6",
   942 => x"1149a275",
   943 => x"cb82c17b",
   944 => x"f304aab7",
   945 => x"c34acc87",
   946 => x"82c17bff",
   947 => x"aab7e0c0",
   948 => x"ff87f404",
   949 => x"78c448d0",
   950 => x"c57bffc3",
   951 => x"7bd3c178",
   952 => x"78c47bc1",
   953 => x"b7c04866",
   954 => x"f0c206a8",
   955 => x"f8e9c287",
   956 => x"66c44cbf",
   957 => x"c8887448",
   958 => x"9c7458a6",
   959 => x"87f9c102",
   960 => x"7efadcc2",
   961 => x"8c4dc0c8",
   962 => x"03acb7c0",
   963 => x"c0c887c6",
   964 => x"4cc04da4",
   965 => x"97ebe9c2",
   966 => x"99d049bf",
   967 => x"c087d102",
   968 => x"f0e9c21e",
   969 => x"87cce849",
   970 => x"497086c4",
   971 => x"87eec04a",
   972 => x"1efadcc2",
   973 => x"49f0e9c2",
   974 => x"c487f9e7",
   975 => x"4a497086",
   976 => x"c848d0ff",
   977 => x"d4c178c5",
   978 => x"bf976e7b",
   979 => x"c1486e7b",
   980 => x"c17e7080",
   981 => x"f0ff058d",
   982 => x"48d0ff87",
   983 => x"9a7278c4",
   984 => x"c087c505",
   985 => x"87c7c148",
   986 => x"e9c21ec1",
   987 => x"e9e549f0",
   988 => x"7486c487",
   989 => x"c7fe059c",
   990 => x"4866c487",
   991 => x"06a8b7c0",
   992 => x"e9c287d1",
   993 => x"78c048f0",
   994 => x"78c080d0",
   995 => x"e9c280f4",
   996 => x"c478bffc",
   997 => x"b7c04866",
   998 => x"d0fd01a8",
   999 => x"48d0ff87",
  1000 => x"d3c178c5",
  1001 => x"c47bc07b",
  1002 => x"c248c178",
  1003 => x"f848c087",
  1004 => x"264d268e",
  1005 => x"264b264c",
  1006 => x"5b5e0e4f",
  1007 => x"1e0e5d5c",
  1008 => x"4cc04b71",
  1009 => x"c004ab4d",
  1010 => x"f7c087e8",
  1011 => x"9d751ed5",
  1012 => x"c087c402",
  1013 => x"c187c24a",
  1014 => x"eb49724a",
  1015 => x"86c487ec",
  1016 => x"84c17e70",
  1017 => x"87c2056e",
  1018 => x"85c14c73",
  1019 => x"ff06ac73",
  1020 => x"486e87d8",
  1021 => x"87f9fe26",
  1022 => x"5c5b5e0e",
  1023 => x"cc4b710e",
  1024 => x"87d80266",
  1025 => x"8cf0c04c",
  1026 => x"7487d802",
  1027 => x"028ac14a",
  1028 => x"028a87d1",
  1029 => x"028a87cd",
  1030 => x"87d987c9",
  1031 => x"e2f94973",
  1032 => x"7487d287",
  1033 => x"c149c01e",
  1034 => x"7487e6d9",
  1035 => x"c149731e",
  1036 => x"c887ded9",
  1037 => x"87fbfd86",
  1038 => x"5c5b5e0e",
  1039 => x"711e0e5d",
  1040 => x"91de494c",
  1041 => x"4dd8eac2",
  1042 => x"6d978571",
  1043 => x"87ddc102",
  1044 => x"bfc4eac2",
  1045 => x"7282744a",
  1046 => x"87ddfd49",
  1047 => x"98487e70",
  1048 => x"87f2c002",
  1049 => x"4bcceac2",
  1050 => x"49cb4a70",
  1051 => x"87f7c0ff",
  1052 => x"93cb4b74",
  1053 => x"83dce5c1",
  1054 => x"c2c183c4",
  1055 => x"49747bf1",
  1056 => x"87f9c2c1",
  1057 => x"e5c17b75",
  1058 => x"49bf97c9",
  1059 => x"cceac21e",
  1060 => x"87e4fd49",
  1061 => x"497486c4",
  1062 => x"87e1c2c1",
  1063 => x"c4c149c0",
  1064 => x"e9c287c0",
  1065 => x"78c048ec",
  1066 => x"dede49c1",
  1067 => x"c0fc2687",
  1068 => x"616f4c87",
  1069 => x"676e6964",
  1070 => x"002e2e2e",
  1071 => x"5c5b5e0e",
  1072 => x"4a4b710e",
  1073 => x"bfc4eac2",
  1074 => x"fb497282",
  1075 => x"4c7087eb",
  1076 => x"87c4029c",
  1077 => x"87fae649",
  1078 => x"48c4eac2",
  1079 => x"49c178c0",
  1080 => x"fb87e8dd",
  1081 => x"5e0e87cd",
  1082 => x"0e5d5c5b",
  1083 => x"dcc286f4",
  1084 => x"4cc04dfa",
  1085 => x"c048a6c4",
  1086 => x"c4eac278",
  1087 => x"a9c049bf",
  1088 => x"87c1c106",
  1089 => x"48fadcc2",
  1090 => x"f8c00298",
  1091 => x"d5f7c087",
  1092 => x"0266c81e",
  1093 => x"a6c487c7",
  1094 => x"c578c048",
  1095 => x"48a6c487",
  1096 => x"66c478c1",
  1097 => x"87e2e649",
  1098 => x"4d7086c4",
  1099 => x"66c484c1",
  1100 => x"c880c148",
  1101 => x"eac258a6",
  1102 => x"ac49bfc4",
  1103 => x"7587c603",
  1104 => x"c8ff059d",
  1105 => x"754cc087",
  1106 => x"e0c3029d",
  1107 => x"d5f7c087",
  1108 => x"0266c81e",
  1109 => x"a6cc87c7",
  1110 => x"c578c048",
  1111 => x"48a6cc87",
  1112 => x"66cc78c1",
  1113 => x"87e2e549",
  1114 => x"7e7086c4",
  1115 => x"c2029848",
  1116 => x"cb4987e8",
  1117 => x"49699781",
  1118 => x"c10299d0",
  1119 => x"c2c187d6",
  1120 => x"49744afc",
  1121 => x"e5c191cb",
  1122 => x"797281dc",
  1123 => x"ffc381c8",
  1124 => x"de497451",
  1125 => x"d8eac291",
  1126 => x"c285714d",
  1127 => x"c17d97c1",
  1128 => x"e0c049a5",
  1129 => x"cae5c251",
  1130 => x"d202bf97",
  1131 => x"c284c187",
  1132 => x"e5c24ba5",
  1133 => x"49db4aca",
  1134 => x"87ebfbfe",
  1135 => x"cd87dbc1",
  1136 => x"51c049a5",
  1137 => x"a5c284c1",
  1138 => x"cb4a6e4b",
  1139 => x"d6fbfe49",
  1140 => x"87c6c187",
  1141 => x"4af8c0c1",
  1142 => x"91cb4974",
  1143 => x"81dce5c1",
  1144 => x"e5c27972",
  1145 => x"02bf97ca",
  1146 => x"497487d8",
  1147 => x"84c191de",
  1148 => x"4bd8eac2",
  1149 => x"e5c28371",
  1150 => x"49dd4aca",
  1151 => x"87e7fafe",
  1152 => x"4b7487d8",
  1153 => x"eac293de",
  1154 => x"a3cb83d8",
  1155 => x"c151c049",
  1156 => x"4a6e7384",
  1157 => x"fafe49cb",
  1158 => x"66c487cd",
  1159 => x"c880c148",
  1160 => x"acc758a6",
  1161 => x"87c5c003",
  1162 => x"e0fc056e",
  1163 => x"f4487487",
  1164 => x"87fdf58e",
  1165 => x"711e731e",
  1166 => x"91cb494b",
  1167 => x"81dce5c1",
  1168 => x"c14aa1c8",
  1169 => x"1248c8e5",
  1170 => x"4aa1c950",
  1171 => x"48c2fac0",
  1172 => x"81ca5012",
  1173 => x"48c9e5c1",
  1174 => x"e5c15011",
  1175 => x"49bf97c9",
  1176 => x"f649c01e",
  1177 => x"e9c287d2",
  1178 => x"78de48ec",
  1179 => x"dad749c1",
  1180 => x"c0f52687",
  1181 => x"4a711e87",
  1182 => x"c191cb49",
  1183 => x"c881dce5",
  1184 => x"c2481181",
  1185 => x"c258f0e9",
  1186 => x"c048c4ea",
  1187 => x"d649c178",
  1188 => x"4f2687f9",
  1189 => x"c049c01e",
  1190 => x"2687c7fc",
  1191 => x"99711e4f",
  1192 => x"c187d202",
  1193 => x"c048f1e6",
  1194 => x"c180f750",
  1195 => x"c140f5c9",
  1196 => x"ce78d5e5",
  1197 => x"ede6c187",
  1198 => x"cee5c148",
  1199 => x"c180fc78",
  1200 => x"2678d4ca",
  1201 => x"5b5e0e4f",
  1202 => x"f40e5d5c",
  1203 => x"494d7186",
  1204 => x"e5c191cb",
  1205 => x"a1c881dc",
  1206 => x"7ea1ca4a",
  1207 => x"c248a6c4",
  1208 => x"78bff4ed",
  1209 => x"4bbf976e",
  1210 => x"734866c4",
  1211 => x"4c4b7028",
  1212 => x"a6cc4812",
  1213 => x"c19c7058",
  1214 => x"9781c984",
  1215 => x"acb74969",
  1216 => x"c087c204",
  1217 => x"bf976e4c",
  1218 => x"4966c84a",
  1219 => x"b9ff3172",
  1220 => x"749966c4",
  1221 => x"70307248",
  1222 => x"b071484a",
  1223 => x"58f8edc2",
  1224 => x"87d9e6c0",
  1225 => x"e2d449c0",
  1226 => x"c0497587",
  1227 => x"f487cef8",
  1228 => x"87fdf18e",
  1229 => x"711e731e",
  1230 => x"c8fe494b",
  1231 => x"fe497387",
  1232 => x"f0f187c3",
  1233 => x"1e731e87",
  1234 => x"a3c64b71",
  1235 => x"87db024a",
  1236 => x"d6028ac1",
  1237 => x"c1028a87",
  1238 => x"028a87da",
  1239 => x"8a87fcc0",
  1240 => x"87e1c002",
  1241 => x"87cb028a",
  1242 => x"c787dbc1",
  1243 => x"87c5fc49",
  1244 => x"c287dec1",
  1245 => x"02bfc4ea",
  1246 => x"4887cbc1",
  1247 => x"eac288c1",
  1248 => x"c1c158c8",
  1249 => x"c8eac287",
  1250 => x"f9c002bf",
  1251 => x"c4eac287",
  1252 => x"80c148bf",
  1253 => x"58c8eac2",
  1254 => x"c287ebc0",
  1255 => x"49bfc4ea",
  1256 => x"eac289c6",
  1257 => x"b7c059c8",
  1258 => x"87da03a9",
  1259 => x"48c4eac2",
  1260 => x"87d278c0",
  1261 => x"bfc8eac2",
  1262 => x"c287cb02",
  1263 => x"48bfc4ea",
  1264 => x"eac280c6",
  1265 => x"49c058c8",
  1266 => x"7387c0d2",
  1267 => x"ecf5c049",
  1268 => x"87e1ef87",
  1269 => x"5c5b5e0e",
  1270 => x"d0ff0e5d",
  1271 => x"59a6dc86",
  1272 => x"c048a6c8",
  1273 => x"c180c478",
  1274 => x"c47866c4",
  1275 => x"c478c180",
  1276 => x"c278c180",
  1277 => x"c148c8ea",
  1278 => x"ece9c278",
  1279 => x"a8de48bf",
  1280 => x"f387cb05",
  1281 => x"497087e0",
  1282 => x"cf59a6cc",
  1283 => x"fde287fc",
  1284 => x"87dfe387",
  1285 => x"7087ece2",
  1286 => x"acfbc04c",
  1287 => x"87fbc102",
  1288 => x"c10566d8",
  1289 => x"c0c187ed",
  1290 => x"82c44a66",
  1291 => x"1e727e6a",
  1292 => x"48ffe0c1",
  1293 => x"c84966c4",
  1294 => x"41204aa1",
  1295 => x"f905aa71",
  1296 => x"26511087",
  1297 => x"66c0c14a",
  1298 => x"f4c8c148",
  1299 => x"c7496a78",
  1300 => x"c1517481",
  1301 => x"c84966c0",
  1302 => x"c151c181",
  1303 => x"c94966c0",
  1304 => x"c151c081",
  1305 => x"ca4966c0",
  1306 => x"c151c081",
  1307 => x"6a1ed81e",
  1308 => x"e281c849",
  1309 => x"86c887d1",
  1310 => x"4866c4c1",
  1311 => x"c701a8c0",
  1312 => x"48a6c887",
  1313 => x"87ce78c1",
  1314 => x"4866c4c1",
  1315 => x"a6d088c1",
  1316 => x"e187c358",
  1317 => x"a6d087dd",
  1318 => x"7478c248",
  1319 => x"e5cd029c",
  1320 => x"4866c887",
  1321 => x"a866c8c1",
  1322 => x"87dacd03",
  1323 => x"c048a6dc",
  1324 => x"c080e878",
  1325 => x"87cbe078",
  1326 => x"d0c14c70",
  1327 => x"dac205ac",
  1328 => x"7e66c487",
  1329 => x"7087efe2",
  1330 => x"59a6c849",
  1331 => x"87f3dfff",
  1332 => x"ecc04c70",
  1333 => x"edc105ac",
  1334 => x"4966c887",
  1335 => x"c0c191cb",
  1336 => x"a1c48166",
  1337 => x"c84d6a4a",
  1338 => x"66c44aa1",
  1339 => x"f5c9c152",
  1340 => x"cedfff79",
  1341 => x"9c4c7087",
  1342 => x"c087d902",
  1343 => x"d302acfb",
  1344 => x"ff557487",
  1345 => x"7087fcde",
  1346 => x"c7029c4c",
  1347 => x"acfbc087",
  1348 => x"87edff05",
  1349 => x"c255e0c0",
  1350 => x"97c055c1",
  1351 => x"4966d87d",
  1352 => x"db05a96e",
  1353 => x"4866c887",
  1354 => x"04a866cc",
  1355 => x"66c887ca",
  1356 => x"cc80c148",
  1357 => x"87c858a6",
  1358 => x"c14866cc",
  1359 => x"58a6d088",
  1360 => x"87ffddff",
  1361 => x"d0c14c70",
  1362 => x"87c805ac",
  1363 => x"c14866d4",
  1364 => x"58a6d880",
  1365 => x"02acd0c1",
  1366 => x"c087e6fd",
  1367 => x"d848a6e0",
  1368 => x"66c47866",
  1369 => x"66e0c048",
  1370 => x"ebc905a8",
  1371 => x"a6e4c087",
  1372 => x"7478c048",
  1373 => x"88fbc048",
  1374 => x"98487e70",
  1375 => x"87edc902",
  1376 => x"7088cb48",
  1377 => x"0298487e",
  1378 => x"4887cdc1",
  1379 => x"7e7088c9",
  1380 => x"c4029848",
  1381 => x"c44887c1",
  1382 => x"487e7088",
  1383 => x"87ce0298",
  1384 => x"7088c148",
  1385 => x"0298487e",
  1386 => x"c887ecc3",
  1387 => x"a6dc87e1",
  1388 => x"78f0c048",
  1389 => x"87cbdcff",
  1390 => x"ecc04c70",
  1391 => x"c4c002ac",
  1392 => x"a6e0c087",
  1393 => x"acecc05c",
  1394 => x"ff87cd02",
  1395 => x"7087f4db",
  1396 => x"acecc04c",
  1397 => x"87f3ff05",
  1398 => x"02acecc0",
  1399 => x"ff87c4c0",
  1400 => x"c087e0db",
  1401 => x"d01eca1e",
  1402 => x"91cb4966",
  1403 => x"4866c8c1",
  1404 => x"a6cc8071",
  1405 => x"4866c858",
  1406 => x"a6d080c4",
  1407 => x"bf66cc58",
  1408 => x"c2dcff49",
  1409 => x"de1ec187",
  1410 => x"bf66d41e",
  1411 => x"f6dbff49",
  1412 => x"7086d087",
  1413 => x"8909c049",
  1414 => x"59a6ecc0",
  1415 => x"4866e8c0",
  1416 => x"c006a8c0",
  1417 => x"e8c087ee",
  1418 => x"a8dd4866",
  1419 => x"87e4c003",
  1420 => x"49bf66c4",
  1421 => x"8166e8c0",
  1422 => x"c051e0c0",
  1423 => x"c14966e8",
  1424 => x"bf66c481",
  1425 => x"51c1c281",
  1426 => x"4966e8c0",
  1427 => x"66c481c2",
  1428 => x"51c081bf",
  1429 => x"c8c1486e",
  1430 => x"496e78f4",
  1431 => x"66d081c8",
  1432 => x"c9496e51",
  1433 => x"5166d481",
  1434 => x"81ca496e",
  1435 => x"d05166dc",
  1436 => x"80c14866",
  1437 => x"c858a6d4",
  1438 => x"66cc4866",
  1439 => x"cbc004a8",
  1440 => x"4866c887",
  1441 => x"a6cc80c1",
  1442 => x"87e1c558",
  1443 => x"c14866cc",
  1444 => x"58a6d088",
  1445 => x"ff87d6c5",
  1446 => x"7087dbdb",
  1447 => x"a6ecc049",
  1448 => x"d1dbff59",
  1449 => x"c0497087",
  1450 => x"dc59a6e0",
  1451 => x"ecc04866",
  1452 => x"cac005a8",
  1453 => x"48a6dc87",
  1454 => x"7866e8c0",
  1455 => x"ff87c4c0",
  1456 => x"c887c0d8",
  1457 => x"91cb4966",
  1458 => x"4866c0c1",
  1459 => x"7e708071",
  1460 => x"6e82c84a",
  1461 => x"c081ca49",
  1462 => x"dc5166e8",
  1463 => x"81c14966",
  1464 => x"8966e8c0",
  1465 => x"307148c1",
  1466 => x"89c14970",
  1467 => x"c27a9771",
  1468 => x"49bff4ed",
  1469 => x"2966e8c0",
  1470 => x"484a6a97",
  1471 => x"f0c09871",
  1472 => x"496e58a6",
  1473 => x"4d6981c4",
  1474 => x"4866e0c0",
  1475 => x"02a866c4",
  1476 => x"c487c8c0",
  1477 => x"78c048a6",
  1478 => x"c487c5c0",
  1479 => x"78c148a6",
  1480 => x"c01e66c4",
  1481 => x"49751ee0",
  1482 => x"87dbd7ff",
  1483 => x"4c7086c8",
  1484 => x"06acb7c0",
  1485 => x"7487d4c1",
  1486 => x"49e0c085",
  1487 => x"4b758974",
  1488 => x"4ac8e1c1",
  1489 => x"dee5fe71",
  1490 => x"c085c287",
  1491 => x"c14866e4",
  1492 => x"a6e8c080",
  1493 => x"66ecc058",
  1494 => x"7081c149",
  1495 => x"c8c002a9",
  1496 => x"48a6c487",
  1497 => x"c5c078c0",
  1498 => x"48a6c487",
  1499 => x"66c478c1",
  1500 => x"49a4c21e",
  1501 => x"7148e0c0",
  1502 => x"1e497088",
  1503 => x"d6ff4975",
  1504 => x"86c887c5",
  1505 => x"01a8b7c0",
  1506 => x"c087c0ff",
  1507 => x"c00266e4",
  1508 => x"496e87d1",
  1509 => x"e4c081c9",
  1510 => x"486e5166",
  1511 => x"78c5cbc1",
  1512 => x"6e87ccc0",
  1513 => x"c281c949",
  1514 => x"c1486e51",
  1515 => x"c878f4cc",
  1516 => x"66cc4866",
  1517 => x"cbc004a8",
  1518 => x"4866c887",
  1519 => x"a6cc80c1",
  1520 => x"87e9c058",
  1521 => x"c14866cc",
  1522 => x"58a6d088",
  1523 => x"ff87dec0",
  1524 => x"7087e0d4",
  1525 => x"87d5c04c",
  1526 => x"05acc6c1",
  1527 => x"d087c8c0",
  1528 => x"80c14866",
  1529 => x"ff58a6d4",
  1530 => x"7087c8d4",
  1531 => x"4866d44c",
  1532 => x"a6d880c1",
  1533 => x"029c7458",
  1534 => x"c887cbc0",
  1535 => x"c8c14866",
  1536 => x"f204a866",
  1537 => x"d3ff87e6",
  1538 => x"66c887e0",
  1539 => x"03a8c748",
  1540 => x"c287e5c0",
  1541 => x"c048c8ea",
  1542 => x"4966c878",
  1543 => x"c0c191cb",
  1544 => x"a1c48166",
  1545 => x"c04a6a4a",
  1546 => x"66c87952",
  1547 => x"cc80c148",
  1548 => x"a8c758a6",
  1549 => x"87dbff04",
  1550 => x"ff8ed0ff",
  1551 => x"4c87f2dd",
  1552 => x"2064616f",
  1553 => x"00202e2a",
  1554 => x"1e00203a",
  1555 => x"4b711e73",
  1556 => x"87c6029b",
  1557 => x"48c4eac2",
  1558 => x"1ec778c0",
  1559 => x"bfc4eac2",
  1560 => x"e5c11e49",
  1561 => x"e9c21edc",
  1562 => x"ed49bfec",
  1563 => x"86cc87e6",
  1564 => x"bfece9c2",
  1565 => x"87e5e849",
  1566 => x"c8029b73",
  1567 => x"dce5c187",
  1568 => x"cae4c049",
  1569 => x"ecdcff87",
  1570 => x"1e731e87",
  1571 => x"e5c14bc0",
  1572 => x"50c048c8",
  1573 => x"bfffe6c1",
  1574 => x"e6d7ff49",
  1575 => x"05987087",
  1576 => x"e2c187c4",
  1577 => x"48734bec",
  1578 => x"87c9dcff",
  1579 => x"204d4f52",
  1580 => x"64616f6c",
  1581 => x"20676e69",
  1582 => x"6c696166",
  1583 => x"1e006465",
  1584 => x"c187e3c7",
  1585 => x"87c3fe49",
  1586 => x"87c3e8fe",
  1587 => x"cd029870",
  1588 => x"fef0fe87",
  1589 => x"02987087",
  1590 => x"4ac187c4",
  1591 => x"4ac087c2",
  1592 => x"ce059a72",
  1593 => x"c11ec087",
  1594 => x"c049cfe4",
  1595 => x"c487d8ef",
  1596 => x"c087fe86",
  1597 => x"dae4c11e",
  1598 => x"caefc049",
  1599 => x"fe1ec087",
  1600 => x"497087c7",
  1601 => x"87ffeec0",
  1602 => x"f887dac3",
  1603 => x"534f268e",
  1604 => x"61662044",
  1605 => x"64656c69",
  1606 => x"6f42002e",
  1607 => x"6e69746f",
  1608 => x"2e2e2e67",
  1609 => x"e6c01e00",
  1610 => x"f2c087e3",
  1611 => x"87f687d3",
  1612 => x"c21e4f26",
  1613 => x"c048c4ea",
  1614 => x"ece9c278",
  1615 => x"fd78c048",
  1616 => x"87e187fd",
  1617 => x"4f2648c0",
  1618 => x"00010000",
  1619 => x"20800000",
  1620 => x"74697845",
  1621 => x"42208000",
  1622 => x"006b6361",
  1623 => x"00001038",
  1624 => x"00002a98",
  1625 => x"38000000",
  1626 => x"b6000010",
  1627 => x"0000002a",
  1628 => x"10380000",
  1629 => x"2ad40000",
  1630 => x"00000000",
  1631 => x"00103800",
  1632 => x"002af200",
  1633 => x"00000000",
  1634 => x"00001038",
  1635 => x"00002b10",
  1636 => x"38000000",
  1637 => x"2e000010",
  1638 => x"0000002b",
  1639 => x"10380000",
  1640 => x"2b4c0000",
  1641 => x"00000000",
  1642 => x"00127500",
  1643 => x"00000000",
  1644 => x"00000000",
  1645 => x"00001345",
  1646 => x"00000000",
  1647 => x"c3000000",
  1648 => x"53000019",
  1649 => x"4944524f",
  1650 => x"5220544e",
  1651 => x"1e004d4f",
  1652 => x"c048f0fe",
  1653 => x"7909cd78",
  1654 => x"1e4f2609",
  1655 => x"bff0fe1e",
  1656 => x"2626487e",
  1657 => x"f0fe1e4f",
  1658 => x"2678c148",
  1659 => x"f0fe1e4f",
  1660 => x"2678c048",
  1661 => x"4a711e4f",
  1662 => x"265252c0",
  1663 => x"5b5e0e4f",
  1664 => x"f40e5d5c",
  1665 => x"974d7186",
  1666 => x"a5c17e6d",
  1667 => x"486c974c",
  1668 => x"6e58a6c8",
  1669 => x"a866c448",
  1670 => x"ff87c505",
  1671 => x"87e6c048",
  1672 => x"c287caff",
  1673 => x"6c9749a5",
  1674 => x"4ba3714b",
  1675 => x"974b6b97",
  1676 => x"486e7e6c",
  1677 => x"a6c880c1",
  1678 => x"cc98c758",
  1679 => x"977058a6",
  1680 => x"87e1fe7c",
  1681 => x"8ef44873",
  1682 => x"4c264d26",
  1683 => x"4f264b26",
  1684 => x"5c5b5e0e",
  1685 => x"7186f40e",
  1686 => x"4a66d84c",
  1687 => x"c29affc3",
  1688 => x"6c974ba4",
  1689 => x"49a17349",
  1690 => x"6c975172",
  1691 => x"c1486e7e",
  1692 => x"58a6c880",
  1693 => x"a6cc98c7",
  1694 => x"f4547058",
  1695 => x"87caff8e",
  1696 => x"e8fd1e1e",
  1697 => x"4abfe087",
  1698 => x"c0e0c049",
  1699 => x"87cb0299",
  1700 => x"edc21e72",
  1701 => x"f7fe49ea",
  1702 => x"fc86c487",
  1703 => x"7e7087fd",
  1704 => x"2687c2fd",
  1705 => x"c21e4f26",
  1706 => x"fd49eaed",
  1707 => x"eac187c7",
  1708 => x"dafc49c0",
  1709 => x"87f7c387",
  1710 => x"5e0e4f26",
  1711 => x"0e5d5c5b",
  1712 => x"edc24d71",
  1713 => x"f4fc49ea",
  1714 => x"c04b7087",
  1715 => x"c304abb7",
  1716 => x"f0c387c2",
  1717 => x"87c905ab",
  1718 => x"48deeec1",
  1719 => x"e3c278c1",
  1720 => x"abe0c387",
  1721 => x"c187c905",
  1722 => x"c148e2ee",
  1723 => x"87d4c278",
  1724 => x"bfe2eec1",
  1725 => x"c287c602",
  1726 => x"c24ca3c0",
  1727 => x"c14c7387",
  1728 => x"02bfdeee",
  1729 => x"7487e0c0",
  1730 => x"29b7c449",
  1731 => x"feefc191",
  1732 => x"cf4a7481",
  1733 => x"c192c29a",
  1734 => x"70307248",
  1735 => x"72baff4a",
  1736 => x"70986948",
  1737 => x"7487db79",
  1738 => x"29b7c449",
  1739 => x"feefc191",
  1740 => x"cf4a7481",
  1741 => x"c392c29a",
  1742 => x"70307248",
  1743 => x"b069484a",
  1744 => x"9d757970",
  1745 => x"87f0c005",
  1746 => x"c848d0ff",
  1747 => x"d4ff78e1",
  1748 => x"c178c548",
  1749 => x"02bfe2ee",
  1750 => x"e0c387c3",
  1751 => x"deeec178",
  1752 => x"87c602bf",
  1753 => x"c348d4ff",
  1754 => x"d4ff78f0",
  1755 => x"ff787348",
  1756 => x"e1c848d0",
  1757 => x"78e0c078",
  1758 => x"48e2eec1",
  1759 => x"eec178c0",
  1760 => x"78c048de",
  1761 => x"49eaedc2",
  1762 => x"7087f2f9",
  1763 => x"abb7c04b",
  1764 => x"87fefc03",
  1765 => x"4d2648c0",
  1766 => x"4b264c26",
  1767 => x"00004f26",
  1768 => x"00000000",
  1769 => x"711e0000",
  1770 => x"cdfc494a",
  1771 => x"1e4f2687",
  1772 => x"49724ac0",
  1773 => x"efc191c4",
  1774 => x"79c081fe",
  1775 => x"b7d082c1",
  1776 => x"87ee04aa",
  1777 => x"5e0e4f26",
  1778 => x"0e5d5c5b",
  1779 => x"dcf84d71",
  1780 => x"c44a7587",
  1781 => x"c1922ab7",
  1782 => x"7582feef",
  1783 => x"c29ccf4c",
  1784 => x"4b496a94",
  1785 => x"9bc32b74",
  1786 => x"307448c2",
  1787 => x"bcff4c70",
  1788 => x"98714874",
  1789 => x"ecf77a70",
  1790 => x"fe487387",
  1791 => x"000087d8",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"00000000",
  1807 => x"ff1e0000",
  1808 => x"e1c848d0",
  1809 => x"ff487178",
  1810 => x"267808d4",
  1811 => x"d0ff1e4f",
  1812 => x"78e1c848",
  1813 => x"d4ff4871",
  1814 => x"66c47808",
  1815 => x"08d4ff48",
  1816 => x"1e4f2678",
  1817 => x"66c44a71",
  1818 => x"49721e49",
  1819 => x"ff87deff",
  1820 => x"e0c048d0",
  1821 => x"4f262678",
  1822 => x"711e731e",
  1823 => x"4966c84b",
  1824 => x"c14a731e",
  1825 => x"ff49a2e0",
  1826 => x"c42687d9",
  1827 => x"264d2687",
  1828 => x"264b264c",
  1829 => x"1e731e4f",
  1830 => x"c24b4a71",
  1831 => x"c803abb7",
  1832 => x"4a49a387",
  1833 => x"c79affc3",
  1834 => x"49a3ce87",
  1835 => x"9affc34a",
  1836 => x"1e4966c8",
  1837 => x"eafe4972",
  1838 => x"d4ff2687",
  1839 => x"d4ff1e87",
  1840 => x"7affc34a",
  1841 => x"c048d0ff",
  1842 => x"7ade78e1",
  1843 => x"bff4edc2",
  1844 => x"c848497a",
  1845 => x"717a7028",
  1846 => x"7028d048",
  1847 => x"d848717a",
  1848 => x"ff7a7028",
  1849 => x"e0c048d0",
  1850 => x"1e4f2678",
  1851 => x"c848d0ff",
  1852 => x"487178c9",
  1853 => x"7808d4ff",
  1854 => x"711e4f26",
  1855 => x"87eb494a",
  1856 => x"c848d0ff",
  1857 => x"1e4f2678",
  1858 => x"4b711e73",
  1859 => x"bfc4eec2",
  1860 => x"c287c302",
  1861 => x"d0ff87eb",
  1862 => x"78c9c848",
  1863 => x"e0c04973",
  1864 => x"48d4ffb1",
  1865 => x"edc27871",
  1866 => x"78c048f8",
  1867 => x"c50266c8",
  1868 => x"49ffc387",
  1869 => x"49c087c2",
  1870 => x"59c0eec2",
  1871 => x"c60266cc",
  1872 => x"d5d5c587",
  1873 => x"cf87c44a",
  1874 => x"c24affff",
  1875 => x"c25ac4ee",
  1876 => x"c148c4ee",
  1877 => x"2687c478",
  1878 => x"264c264d",
  1879 => x"0e4f264b",
  1880 => x"5d5c5b5e",
  1881 => x"c24a710e",
  1882 => x"4cbfc0ee",
  1883 => x"cb029a72",
  1884 => x"91c84987",
  1885 => x"4bfdf3c1",
  1886 => x"87c48371",
  1887 => x"4bfdf7c1",
  1888 => x"49134dc0",
  1889 => x"edc29974",
  1890 => x"ffb9bffc",
  1891 => x"787148d4",
  1892 => x"852cb7c1",
  1893 => x"04adb7c8",
  1894 => x"edc287e8",
  1895 => x"c848bff8",
  1896 => x"fcedc280",
  1897 => x"87effe58",
  1898 => x"711e731e",
  1899 => x"9a4a134b",
  1900 => x"7287cb02",
  1901 => x"87e7fe49",
  1902 => x"059a4a13",
  1903 => x"dafe87f5",
  1904 => x"edc21e87",
  1905 => x"c249bff8",
  1906 => x"c148f8ed",
  1907 => x"c0c478a1",
  1908 => x"db03a9b7",
  1909 => x"48d4ff87",
  1910 => x"bffcedc2",
  1911 => x"f8edc278",
  1912 => x"edc249bf",
  1913 => x"a1c148f8",
  1914 => x"b7c0c478",
  1915 => x"87e504a9",
  1916 => x"c848d0ff",
  1917 => x"c4eec278",
  1918 => x"2678c048",
  1919 => x"0000004f",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00005f5f",
  1923 => x"03030000",
  1924 => x"00030300",
  1925 => x"7f7f1400",
  1926 => x"147f7f14",
  1927 => x"2e240000",
  1928 => x"123a6b6b",
  1929 => x"366a4c00",
  1930 => x"32566c18",
  1931 => x"4f7e3000",
  1932 => x"683a7759",
  1933 => x"04000040",
  1934 => x"00000307",
  1935 => x"1c000000",
  1936 => x"0041633e",
  1937 => x"41000000",
  1938 => x"001c3e63",
  1939 => x"3e2a0800",
  1940 => x"2a3e1c1c",
  1941 => x"08080008",
  1942 => x"08083e3e",
  1943 => x"80000000",
  1944 => x"000060e0",
  1945 => x"08080000",
  1946 => x"08080808",
  1947 => x"00000000",
  1948 => x"00006060",
  1949 => x"30604000",
  1950 => x"03060c18",
  1951 => x"7f3e0001",
  1952 => x"3e7f4d59",
  1953 => x"06040000",
  1954 => x"00007f7f",
  1955 => x"63420000",
  1956 => x"464f5971",
  1957 => x"63220000",
  1958 => x"367f4949",
  1959 => x"161c1800",
  1960 => x"107f7f13",
  1961 => x"67270000",
  1962 => x"397d4545",
  1963 => x"7e3c0000",
  1964 => x"3079494b",
  1965 => x"01010000",
  1966 => x"070f7971",
  1967 => x"7f360000",
  1968 => x"367f4949",
  1969 => x"4f060000",
  1970 => x"1e3f6949",
  1971 => x"00000000",
  1972 => x"00006666",
  1973 => x"80000000",
  1974 => x"000066e6",
  1975 => x"08080000",
  1976 => x"22221414",
  1977 => x"14140000",
  1978 => x"14141414",
  1979 => x"22220000",
  1980 => x"08081414",
  1981 => x"03020000",
  1982 => x"060f5951",
  1983 => x"417f3e00",
  1984 => x"1e1f555d",
  1985 => x"7f7e0000",
  1986 => x"7e7f0909",
  1987 => x"7f7f0000",
  1988 => x"367f4949",
  1989 => x"3e1c0000",
  1990 => x"41414163",
  1991 => x"7f7f0000",
  1992 => x"1c3e6341",
  1993 => x"7f7f0000",
  1994 => x"41414949",
  1995 => x"7f7f0000",
  1996 => x"01010909",
  1997 => x"7f3e0000",
  1998 => x"7a7b4941",
  1999 => x"7f7f0000",
  2000 => x"7f7f0808",
  2001 => x"41000000",
  2002 => x"00417f7f",
  2003 => x"60200000",
  2004 => x"3f7f4040",
  2005 => x"087f7f00",
  2006 => x"4163361c",
  2007 => x"7f7f0000",
  2008 => x"40404040",
  2009 => x"067f7f00",
  2010 => x"7f7f060c",
  2011 => x"067f7f00",
  2012 => x"7f7f180c",
  2013 => x"7f3e0000",
  2014 => x"3e7f4141",
  2015 => x"7f7f0000",
  2016 => x"060f0909",
  2017 => x"417f3e00",
  2018 => x"407e7f61",
  2019 => x"7f7f0000",
  2020 => x"667f1909",
  2021 => x"6f260000",
  2022 => x"327b594d",
  2023 => x"01010000",
  2024 => x"01017f7f",
  2025 => x"7f3f0000",
  2026 => x"3f7f4040",
  2027 => x"3f0f0000",
  2028 => x"0f3f7070",
  2029 => x"307f7f00",
  2030 => x"7f7f3018",
  2031 => x"36634100",
  2032 => x"63361c1c",
  2033 => x"06030141",
  2034 => x"03067c7c",
  2035 => x"59716101",
  2036 => x"4143474d",
  2037 => x"7f000000",
  2038 => x"0041417f",
  2039 => x"06030100",
  2040 => x"6030180c",
  2041 => x"41000040",
  2042 => x"007f7f41",
  2043 => x"060c0800",
  2044 => x"080c0603",
  2045 => x"80808000",
  2046 => x"80808080",
  2047 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
