library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"00040703",
     1 => x"74200000",
     2 => x"787c5454",
     3 => x"7f7f0000",
     4 => x"387c4444",
     5 => x"7c380000",
     6 => x"00444444",
     7 => x"7c380000",
     8 => x"7f7f4444",
     9 => x"7c380000",
    10 => x"185c5454",
    11 => x"7e040000",
    12 => x"0005057f",
    13 => x"bc180000",
    14 => x"7cfca4a4",
    15 => x"7f7f0000",
    16 => x"787c0404",
    17 => x"00000000",
    18 => x"00407d3d",
    19 => x"80800000",
    20 => x"007dfd80",
    21 => x"7f7f0000",
    22 => x"446c3810",
    23 => x"00000000",
    24 => x"00407f3f",
    25 => x"0c7c7c00",
    26 => x"787c0c18",
    27 => x"7c7c0000",
    28 => x"787c0404",
    29 => x"7c380000",
    30 => x"387c4444",
    31 => x"fcfc0000",
    32 => x"183c2424",
    33 => x"3c180000",
    34 => x"fcfc2424",
    35 => x"7c7c0000",
    36 => x"080c0404",
    37 => x"5c480000",
    38 => x"20745454",
    39 => x"3f040000",
    40 => x"0044447f",
    41 => x"7c3c0000",
    42 => x"7c7c4040",
    43 => x"3c1c0000",
    44 => x"1c3c6060",
    45 => x"607c3c00",
    46 => x"3c7c6030",
    47 => x"386c4400",
    48 => x"446c3810",
    49 => x"bc1c0000",
    50 => x"1c3c60e0",
    51 => x"64440000",
    52 => x"444c5c74",
    53 => x"08080000",
    54 => x"4141773e",
    55 => x"00000000",
    56 => x"00007f7f",
    57 => x"41410000",
    58 => x"08083e77",
    59 => x"01010200",
    60 => x"01020203",
    61 => x"7f7f7f00",
    62 => x"7f7f7f7f",
    63 => x"1c080800",
    64 => x"7f3e3e1c",
    65 => x"3e7f7f7f",
    66 => x"081c1c3e",
    67 => x"18100008",
    68 => x"10187c7c",
    69 => x"30100000",
    70 => x"10307c7c",
    71 => x"60301000",
    72 => x"061e7860",
    73 => x"3c664200",
    74 => x"42663c18",
    75 => x"6a387800",
    76 => x"386cc6c2",
    77 => x"00006000",
    78 => x"60000060",
    79 => x"5b5e0e00",
    80 => x"1e0e5d5c",
    81 => x"eec24c71",
    82 => x"c04dbfd5",
    83 => x"741ec04b",
    84 => x"87c702ab",
    85 => x"c048a6c4",
    86 => x"c487c578",
    87 => x"78c148a6",
    88 => x"731e66c4",
    89 => x"87dfee49",
    90 => x"e0c086c8",
    91 => x"87efef49",
    92 => x"6a4aa5c4",
    93 => x"87f0f049",
    94 => x"cb87c6f1",
    95 => x"c883c185",
    96 => x"ff04abb7",
    97 => x"262687c7",
    98 => x"264c264d",
    99 => x"1e4f264b",
   100 => x"eec24a71",
   101 => x"eec25ad9",
   102 => x"78c748d9",
   103 => x"87ddfe49",
   104 => x"731e4f26",
   105 => x"c04a711e",
   106 => x"d303aab7",
   107 => x"e0d4c287",
   108 => x"87c405bf",
   109 => x"87c24bc1",
   110 => x"d4c24bc0",
   111 => x"87c45be4",
   112 => x"5ae4d4c2",
   113 => x"bfe0d4c2",
   114 => x"c19ac14a",
   115 => x"ec49a2c0",
   116 => x"48fc87e8",
   117 => x"bfe0d4c2",
   118 => x"87effe78",
   119 => x"c44a711e",
   120 => x"49721e66",
   121 => x"2687eeea",
   122 => x"711e4f26",
   123 => x"48d4ff4a",
   124 => x"ff78ffc3",
   125 => x"e1c048d0",
   126 => x"48d4ff78",
   127 => x"497278c1",
   128 => x"787131c4",
   129 => x"c048d0ff",
   130 => x"4f2678e0",
   131 => x"e0d4c21e",
   132 => x"d1e649bf",
   133 => x"cdeec287",
   134 => x"78bfe848",
   135 => x"48c9eec2",
   136 => x"c278bfec",
   137 => x"4abfcdee",
   138 => x"99ffc349",
   139 => x"722ab7c8",
   140 => x"c2b07148",
   141 => x"2658d5ee",
   142 => x"5b5e0e4f",
   143 => x"710e5d5c",
   144 => x"87c8ff4b",
   145 => x"48c8eec2",
   146 => x"497350c0",
   147 => x"7087f7e5",
   148 => x"9cc24c49",
   149 => x"cb49eecb",
   150 => x"497087ce",
   151 => x"c8eec24d",
   152 => x"c105bf97",
   153 => x"66d087e2",
   154 => x"d1eec249",
   155 => x"d60599bf",
   156 => x"4966d487",
   157 => x"bfc9eec2",
   158 => x"87cb0599",
   159 => x"c5e54973",
   160 => x"02987087",
   161 => x"c187c1c1",
   162 => x"87c0fe4c",
   163 => x"e3ca4975",
   164 => x"02987087",
   165 => x"eec287c6",
   166 => x"50c148c8",
   167 => x"97c8eec2",
   168 => x"e3c005bf",
   169 => x"d1eec287",
   170 => x"66d049bf",
   171 => x"d6ff0599",
   172 => x"c9eec287",
   173 => x"66d449bf",
   174 => x"caff0599",
   175 => x"e4497387",
   176 => x"987087c4",
   177 => x"87fffe05",
   178 => x"fafa4874",
   179 => x"5b5e0e87",
   180 => x"f80e5d5c",
   181 => x"4c4dc086",
   182 => x"c47ebfec",
   183 => x"eec248a6",
   184 => x"c178bfd5",
   185 => x"c71ec01e",
   186 => x"87cdfd49",
   187 => x"987086c8",
   188 => x"ff87cd02",
   189 => x"87eafa49",
   190 => x"e349dac1",
   191 => x"4dc187c8",
   192 => x"97c8eec2",
   193 => x"87cf02bf",
   194 => x"bfd8d4c2",
   195 => x"c2b9c149",
   196 => x"7159dcd4",
   197 => x"c287d3fb",
   198 => x"4bbfcdee",
   199 => x"bfe0d4c2",
   200 => x"87e9c005",
   201 => x"e249fdc3",
   202 => x"fac387dc",
   203 => x"87d6e249",
   204 => x"ffc34973",
   205 => x"c01e7199",
   206 => x"87e0fa49",
   207 => x"b7c84973",
   208 => x"c11e7129",
   209 => x"87d4fa49",
   210 => x"f5c586c8",
   211 => x"d1eec287",
   212 => x"029b4bbf",
   213 => x"d4c287dd",
   214 => x"c749bfdc",
   215 => x"987087d6",
   216 => x"c087c405",
   217 => x"c287d24b",
   218 => x"fbc649e0",
   219 => x"e0d4c287",
   220 => x"c287c658",
   221 => x"c048dcd4",
   222 => x"c2497378",
   223 => x"87cd0599",
   224 => x"e149ebc3",
   225 => x"497087c0",
   226 => x"c20299c2",
   227 => x"734cfb87",
   228 => x"0599c149",
   229 => x"f4c387cd",
   230 => x"87eae049",
   231 => x"99c24970",
   232 => x"fa87c202",
   233 => x"c849734c",
   234 => x"87cd0599",
   235 => x"e049f5c3",
   236 => x"497087d4",
   237 => x"d50299c2",
   238 => x"d9eec287",
   239 => x"87ca02bf",
   240 => x"c288c148",
   241 => x"c058ddee",
   242 => x"4cff87c2",
   243 => x"49734dc1",
   244 => x"ce0599c4",
   245 => x"49f2c387",
   246 => x"87eadfff",
   247 => x"99c24970",
   248 => x"c287dc02",
   249 => x"7ebfd9ee",
   250 => x"a8b7c748",
   251 => x"87cbc003",
   252 => x"80c1486e",
   253 => x"58ddeec2",
   254 => x"fe87c2c0",
   255 => x"c34dc14c",
   256 => x"dfff49fd",
   257 => x"497087c0",
   258 => x"d50299c2",
   259 => x"d9eec287",
   260 => x"c9c002bf",
   261 => x"d9eec287",
   262 => x"c078c048",
   263 => x"4cfd87c2",
   264 => x"fac34dc1",
   265 => x"dddeff49",
   266 => x"c2497087",
   267 => x"d9c00299",
   268 => x"d9eec287",
   269 => x"b7c748bf",
   270 => x"c9c003a8",
   271 => x"d9eec287",
   272 => x"c078c748",
   273 => x"4cfc87c2",
   274 => x"b7c04dc1",
   275 => x"d3c003ac",
   276 => x"4866c487",
   277 => x"7080d8c1",
   278 => x"02bf6e7e",
   279 => x"4b87c5c0",
   280 => x"0f734974",
   281 => x"f0c31ec0",
   282 => x"49dac11e",
   283 => x"c887caf7",
   284 => x"02987086",
   285 => x"c287d8c0",
   286 => x"7ebfd9ee",
   287 => x"91cb496e",
   288 => x"714a66c4",
   289 => x"c0026a82",
   290 => x"6e4b87c5",
   291 => x"750f7349",
   292 => x"c8c0029d",
   293 => x"d9eec287",
   294 => x"e0f249bf",
   295 => x"e4d4c287",
   296 => x"ddc002bf",
   297 => x"cbc24987",
   298 => x"02987087",
   299 => x"c287d3c0",
   300 => x"49bfd9ee",
   301 => x"c087c6f2",
   302 => x"87e6f349",
   303 => x"48e4d4c2",
   304 => x"8ef878c0",
   305 => x"0e87c0f3",
   306 => x"5d5c5b5e",
   307 => x"4c711e0e",
   308 => x"bfd5eec2",
   309 => x"a1cdc149",
   310 => x"81d1c14d",
   311 => x"9c747e69",
   312 => x"c487cf02",
   313 => x"7b744ba5",
   314 => x"bfd5eec2",
   315 => x"87dff249",
   316 => x"9c747b6e",
   317 => x"c087c405",
   318 => x"c187c24b",
   319 => x"f249734b",
   320 => x"66d487e0",
   321 => x"4987c702",
   322 => x"4a7087de",
   323 => x"4ac087c2",
   324 => x"5ae8d4c2",
   325 => x"87eff126",
   326 => x"00000000",
   327 => x"00000000",
   328 => x"00000000",
   329 => x"00000000",
   330 => x"ff4a711e",
   331 => x"7249bfc8",
   332 => x"4f2648a1",
   333 => x"bfc8ff1e",
   334 => x"c0c0fe89",
   335 => x"a9c0c0c0",
   336 => x"c087c401",
   337 => x"c187c24a",
   338 => x"2648724a",
   339 => x"5b5e0e4f",
   340 => x"710e5d5c",
   341 => x"4cd4ff4b",
   342 => x"c04866d0",
   343 => x"ff49d678",
   344 => x"c387dbdb",
   345 => x"496c7cff",
   346 => x"7199ffc3",
   347 => x"f0c3494d",
   348 => x"a9e0c199",
   349 => x"c387cb05",
   350 => x"486c7cff",
   351 => x"66d098c3",
   352 => x"ffc37808",
   353 => x"494a6c7c",
   354 => x"ffc331c8",
   355 => x"714a6c7c",
   356 => x"c84972b2",
   357 => x"7cffc331",
   358 => x"b2714a6c",
   359 => x"31c84972",
   360 => x"6c7cffc3",
   361 => x"ffb2714a",
   362 => x"e0c048d0",
   363 => x"029b7378",
   364 => x"7b7287c2",
   365 => x"4d264875",
   366 => x"4b264c26",
   367 => x"261e4f26",
   368 => x"5b5e0e4f",
   369 => x"86f80e5c",
   370 => x"a6c81e76",
   371 => x"87fdfd49",
   372 => x"4b7086c4",
   373 => x"a8c2486e",
   374 => x"87f0c203",
   375 => x"f0c34a73",
   376 => x"aad0c19a",
   377 => x"c187c702",
   378 => x"c205aae0",
   379 => x"497387de",
   380 => x"c30299c8",
   381 => x"87c6ff87",
   382 => x"9cc34c73",
   383 => x"c105acc2",
   384 => x"66c487c2",
   385 => x"7131c949",
   386 => x"4a66c41e",
   387 => x"eec292d4",
   388 => x"817249dd",
   389 => x"87facefe",
   390 => x"d8ff49d8",
   391 => x"c0c887e0",
   392 => x"fadcc21e",
   393 => x"f5eafd49",
   394 => x"48d0ff87",
   395 => x"c278e0c0",
   396 => x"cc1efadc",
   397 => x"92d44a66",
   398 => x"49ddeec2",
   399 => x"cdfe8172",
   400 => x"86cc87c1",
   401 => x"c105acc1",
   402 => x"66c487c2",
   403 => x"7131c949",
   404 => x"4a66c41e",
   405 => x"eec292d4",
   406 => x"817249dd",
   407 => x"87f2cdfe",
   408 => x"1efadcc2",
   409 => x"d44a66c8",
   410 => x"ddeec292",
   411 => x"fe817249",
   412 => x"d787c1cb",
   413 => x"c5d7ff49",
   414 => x"1ec0c887",
   415 => x"49fadcc2",
   416 => x"87f3e8fd",
   417 => x"d0ff86cc",
   418 => x"78e0c048",
   419 => x"e7fc8ef8",
   420 => x"5b5e0e87",
   421 => x"1e0e5d5c",
   422 => x"d4ff4d71",
   423 => x"7e66d44c",
   424 => x"a8b7c348",
   425 => x"c087c506",
   426 => x"87e2c148",
   427 => x"dbfe4975",
   428 => x"1e7587ed",
   429 => x"d44b66c4",
   430 => x"ddeec293",
   431 => x"fe497383",
   432 => x"c887fdc4",
   433 => x"ff4b6b83",
   434 => x"e1c848d0",
   435 => x"737cdd78",
   436 => x"99ffc349",
   437 => x"49737c71",
   438 => x"c329b7c8",
   439 => x"7c7199ff",
   440 => x"b7d04973",
   441 => x"99ffc329",
   442 => x"49737c71",
   443 => x"7129b7d8",
   444 => x"7c7cc07c",
   445 => x"7c7c7c7c",
   446 => x"7c7c7c7c",
   447 => x"e0c07c7c",
   448 => x"1e66c478",
   449 => x"d5ff49dc",
   450 => x"86c887d9",
   451 => x"fa264873",
   452 => x"fa2687e4",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
